module IFetch(
  input         reset,
  input         io_jump_en,
  input  [63:0] io_jump_pc,
  input  [63:0] io_pc,
  output [63:0] io_next_pc,
  output        io_valid
);
  wire [63:0] _io_next_pc_T_1 = io_pc + 64'h4; // @[IFetch.scala 13:51]
  assign io_next_pc = io_jump_en ? io_jump_pc : _io_next_pc_T_1; // @[IFetch.scala 13:20]
  assign io_valid = ~reset; // @[IFetch.scala 14:17]
endmodule
module Decode(
  input  [63:0] io_pc,
  input  [31:0] io_inst,
  output        io_rs1_en,
  output        io_rs2_en,
  output [4:0]  io_rs1_addr,
  output [4:0]  io_rs2_addr,
  input  [63:0] io_rs1_data,
  input  [63:0] io_rs2_data,
  output        io_rd_en,
  output [4:0]  io_rd_addr,
  output [6:0]  io_decode_info_fu_code,
  output [15:0] io_decode_info_alu_code,
  output [7:0]  io_decode_info_bu_code,
  output [6:0]  io_decode_info_lu_code,
  output [3:0]  io_decode_info_su_code,
  output [1:0]  io_decode_info_mu_code,
  output [7:0]  io_decode_info_du_code,
  output [7:0]  io_decode_info_csru_code,
  output        io_jump_en,
  output [63:0] io_jump_pc,
  output [63:0] io_op1,
  output [63:0] io_op2,
  output [63:0] io_imm,
  output        io_putch,
  input  [63:0] io_mtvec,
  input  [63:0] io_mepc
);
  wire [31:0] _sll_T = io_inst & 32'hfe00707f; // @[Decode.scala 56:20]
  wire  sll = 32'h1033 == _sll_T; // @[Decode.scala 56:20]
  wire  srl = 32'h5033 == _sll_T; // @[Decode.scala 57:20]
  wire  sra = 32'h40005033 == _sll_T; // @[Decode.scala 58:20]
  wire [31:0] _slli_T = io_inst & 32'hfc00707f; // @[Decode.scala 59:21]
  wire  slli = 32'h1013 == _slli_T; // @[Decode.scala 59:21]
  wire  srli = 32'h5013 == _slli_T; // @[Decode.scala 60:21]
  wire  srai = 32'h40005013 == _slli_T; // @[Decode.scala 61:21]
  wire  sllw = 32'h103b == _sll_T; // @[Decode.scala 62:21]
  wire  srlw = 32'h503b == _sll_T; // @[Decode.scala 63:21]
  wire  sraw = 32'h4000503b == _sll_T; // @[Decode.scala 64:21]
  wire  slliw = 32'h101b == _sll_T; // @[Decode.scala 65:22]
  wire  srliw = 32'h501b == _sll_T; // @[Decode.scala 66:22]
  wire  sraiw = 32'h4000501b == _sll_T; // @[Decode.scala 67:22]
  wire  add = 32'h33 == _sll_T; // @[Decode.scala 69:24]
  wire  addw = 32'h3b == _sll_T; // @[Decode.scala 70:24]
  wire [31:0] _addi_T = io_inst & 32'h707f; // @[Decode.scala 71:24]
  wire  addi = 32'h13 == _addi_T; // @[Decode.scala 71:24]
  wire  addiw = 32'h1b == _addi_T; // @[Decode.scala 72:24]
  wire  alu_sub = 32'h40000033 == _sll_T; // @[Decode.scala 73:24]
  wire  alu_subw = 32'h4000003b == _sll_T; // @[Decode.scala 74:24]
  wire [31:0] _lui_T = io_inst & 32'h7f; // @[Decode.scala 75:24]
  wire  lui = 32'h37 == _lui_T; // @[Decode.scala 75:24]
  wire  alu_auipc = 32'h17 == _lui_T; // @[Decode.scala 76:24]
  wire  xor_ = 32'h4033 == _sll_T; // @[Decode.scala 78:24]
  wire  or_ = 32'h6033 == _sll_T; // @[Decode.scala 79:24]
  wire  and_ = 32'h7033 == _sll_T; // @[Decode.scala 80:24]
  wire  xori = 32'h4013 == _addi_T; // @[Decode.scala 81:24]
  wire  ori = 32'h6013 == _addi_T; // @[Decode.scala 82:24]
  wire  andi = 32'h7013 == _addi_T; // @[Decode.scala 83:24]
  wire  slt = 32'h2033 == _sll_T; // @[Decode.scala 85:24]
  wire  sltu = 32'h3033 == _sll_T; // @[Decode.scala 86:24]
  wire  slti = 32'h2013 == _addi_T; // @[Decode.scala 87:24]
  wire  sltiu = 32'h3013 == _addi_T; // @[Decode.scala 88:24]
  wire  beq = 32'h63 == _addi_T; // @[Decode.scala 90:24]
  wire  bne = 32'h1063 == _addi_T; // @[Decode.scala 91:24]
  wire  blt = 32'h4063 == _addi_T; // @[Decode.scala 92:24]
  wire  bge = 32'h5063 == _addi_T; // @[Decode.scala 93:24]
  wire  bltu = 32'h6063 == _addi_T; // @[Decode.scala 94:24]
  wire  bgeu = 32'h7063 == _addi_T; // @[Decode.scala 95:24]
  wire  jal = 32'h6f == _lui_T; // @[Decode.scala 97:24]
  wire  jalr = 32'h67 == _addi_T; // @[Decode.scala 98:24]
  wire  lb = 32'h3 == _addi_T; // @[Decode.scala 100:24]
  wire  lh = 32'h1003 == _addi_T; // @[Decode.scala 101:24]
  wire  lw = 32'h2003 == _addi_T; // @[Decode.scala 102:24]
  wire  ld = 32'h3003 == _addi_T; // @[Decode.scala 103:24]
  wire  lbu = 32'h4003 == _addi_T; // @[Decode.scala 104:24]
  wire  lhu = 32'h5003 == _addi_T; // @[Decode.scala 105:24]
  wire  lwu = 32'h6003 == _addi_T; // @[Decode.scala 106:24]
  wire  sb = 32'h23 == _addi_T; // @[Decode.scala 108:24]
  wire  sh = 32'h1023 == _addi_T; // @[Decode.scala 109:24]
  wire  sw = 32'h2023 == _addi_T; // @[Decode.scala 110:24]
  wire  sd = 32'h3023 == _addi_T; // @[Decode.scala 111:24]
  wire  mul = 32'h2000033 == _sll_T; // @[Decode.scala 113:24]
  wire  mulw = 32'h200003b == _sll_T; // @[Decode.scala 114:24]
  wire  div = 32'h2004033 == _sll_T; // @[Decode.scala 115:24]
  wire  divw = 32'h200403b == _sll_T; // @[Decode.scala 116:24]
  wire  divu = 32'h2005033 == _sll_T; // @[Decode.scala 117:24]
  wire  divuw = 32'h200503b == _sll_T; // @[Decode.scala 118:24]
  wire  rem = 32'h2006033 == _sll_T; // @[Decode.scala 119:24]
  wire  remw = 32'h200603b == _sll_T; // @[Decode.scala 120:24]
  wire  remu = 32'h2007033 == _sll_T; // @[Decode.scala 121:24]
  wire  remuw = 32'h200703b == _sll_T; // @[Decode.scala 122:24]
  wire  ecall = 32'h73 == io_inst; // @[Decode.scala 124:24]
  wire  mret = 32'h30200073 == io_inst; // @[Decode.scala 125:24]
  wire  csrrs = 32'h2073 == _addi_T; // @[Decode.scala 126:24]
  wire  csrrw = 32'h1073 == _addi_T; // @[Decode.scala 127:24]
  wire  csrrc = 32'h3073 == _addi_T; // @[Decode.scala 128:24]
  wire  csrrsi = 32'h6073 == _addi_T; // @[Decode.scala 129:24]
  wire  csrrwi = 32'h5073 == _addi_T; // @[Decode.scala 130:24]
  wire  csrrci = 32'h7073 == _addi_T; // @[Decode.scala 131:24]
  wire  alu_add = add | addi | lui; // @[Decode.scala 139:33]
  wire  alu_addw = addw | addiw; // @[Decode.scala 140:26]
  wire  alu_sll = sll | slli; // @[Decode.scala 145:26]
  wire  alu_srl = srl | srli; // @[Decode.scala 146:26]
  wire  alu_sra = sra | srai; // @[Decode.scala 147:26]
  wire  alu_sllw = sllw | slliw; // @[Decode.scala 148:26]
  wire  alu_srlw = srlw | srliw; // @[Decode.scala 149:26]
  wire  alu_sraw = sraw | sraiw; // @[Decode.scala 150:26]
  wire  alu_xor = xor_ | xori; // @[Decode.scala 152:26]
  wire  alu_or = or_ | ori; // @[Decode.scala 153:26]
  wire  alu_and = and_ | andi; // @[Decode.scala 154:26]
  wire  alu_slt = slt | slti; // @[Decode.scala 156:26]
  wire  alu_sltu = sltu | sltiu; // @[Decode.scala 157:26]
  wire [7:0] alu_code_lo = {alu_sra,alu_srl,alu_sll,alu_auipc,alu_subw,alu_sub,alu_addw,alu_add}; // @[Cat.scala 30:58]
  wire [7:0] alu_code_hi = {alu_sltu,alu_slt,alu_and,alu_or,alu_xor,alu_sraw,alu_srlw,alu_sllw}; // @[Cat.scala 30:58]
  wire [15:0] alu_code = {alu_sltu,alu_slt,alu_and,alu_or,alu_xor,alu_sraw,alu_srlw,alu_sllw,alu_code_lo}; // @[Cat.scala 30:58]
  wire  alu_en = alu_code != 16'h0; // @[Decode.scala 160:29]
  wire [3:0] bu_code_lo = {bge,blt,bne,beq}; // @[Cat.scala 30:58]
  wire [3:0] bu_code_hi = {jalr,jal,bgeu,bltu}; // @[Cat.scala 30:58]
  wire [7:0] bu_code = {jalr,jal,bgeu,bltu,bge,blt,bne,beq}; // @[Cat.scala 30:58]
  wire  bu_en = bu_code != 8'h0; // @[Decode.scala 163:27]
  wire [2:0] lu_code_lo = {lw,lh,lb}; // @[Cat.scala 30:58]
  wire [3:0] lu_code_hi = {lwu,lhu,lbu,ld}; // @[Cat.scala 30:58]
  wire [6:0] lu_code = {lwu,lhu,lbu,ld,lw,lh,lb}; // @[Cat.scala 30:58]
  wire  lu_en = lu_code != 7'h0; // @[Decode.scala 166:27]
  wire [1:0] su_code_lo = {sh,sb}; // @[Cat.scala 30:58]
  wire [1:0] su_code_hi = {sd,sw}; // @[Cat.scala 30:58]
  wire [3:0] su_code = {sd,sw,sh,sb}; // @[Cat.scala 30:58]
  wire  su_en = su_code != 4'h0; // @[Decode.scala 169:27]
  wire [1:0] mu_code = {mulw,mul}; // @[Cat.scala 30:58]
  wire  mu_en = mu_code != 2'h0; // @[Decode.scala 172:27]
  wire [3:0] du_code_lo = {divuw,divu,divw,div}; // @[Cat.scala 30:58]
  wire [3:0] du_code_hi = {remuw,remu,remw,rem}; // @[Cat.scala 30:58]
  wire [7:0] du_code = {remuw,remu,remw,rem,divuw,divu,divw,div}; // @[Cat.scala 30:58]
  wire  du_en = du_code != 8'h0; // @[Decode.scala 175:27]
  wire [3:0] csru_code_lo = {csrrw,csrrs,mret,ecall}; // @[Cat.scala 30:58]
  wire [3:0] csru_code_hi = {csrrci,csrrwi,csrrsi,csrrc}; // @[Cat.scala 30:58]
  wire [7:0] csru_code = {csrrci,csrrwi,csrrsi,csrrc,csrrw,csrrs,mret,ecall}; // @[Cat.scala 30:58]
  wire  csr_en = csru_code != 8'h0; // @[Decode.scala 178:31]
  wire [2:0] fu_code_lo = {lu_en,bu_en,alu_en}; // @[Cat.scala 30:58]
  wire [3:0] fu_code_hi = {csr_en,du_en,mu_en,su_en}; // @[Cat.scala 30:58]
  wire  _type_r_T_5 = sll | srl | sra | sllw | srlw | sraw | add; // @[Decode.scala 183:74]
  wire  _type_r_T_9 = _type_r_T_5 | addw | alu_sub | alu_subw | xor_; // @[Decode.scala 184:54]
  wire  _type_r_T_12 = _type_r_T_9 | or_ | and_ | slt; // @[Decode.scala 185:45]
  wire  _type_r_T_14 = _type_r_T_12 | sltu | mul; // @[Decode.scala 186:36]
  wire  _type_r_T_16 = _type_r_T_14 | mulw | div; // @[Decode.scala 187:36]
  wire  _type_r_T_20 = _type_r_T_16 | divw | divu | divuw | rem; // @[Decode.scala 188:54]
  wire  type_r = _type_r_T_20 | remw | remu | remuw | mret; // @[Decode.scala 189:54]
  wire  _type_i_T_5 = slli | srli | srai | slliw | srliw | sraiw | addi; // @[Decode.scala 191:74]
  wire  _type_i_T_7 = _type_i_T_5 | addiw | xori; // @[Decode.scala 192:36]
  wire  _type_i_T_10 = _type_i_T_7 | ori | andi | slti; // @[Decode.scala 193:45]
  wire  _type_i_T_12 = _type_i_T_10 | sltiu | jalr; // @[Decode.scala 194:36]
  wire  _type_i_T_13 = _type_i_T_12 | lb; // @[Decode.scala 195:27]
  wire  _type_i_T_20 = _type_i_T_13 | lh | lw | ld | lbu | lhu | lwu | ecall; // @[Decode.scala 196:81]
  wire  type_i = _type_i_T_20 | csrrs | csrrw | csrrc | csrrwi | csrrci | csrrsi; // @[Decode.scala 197:74]
  wire  type_s = sb | sh | sw | sd; // @[Decode.scala 198:45]
  wire  type_b = beq | bne | blt | bge | bltu | bgeu; // @[Decode.scala 199:64]
  wire  type_u = lui | alu_auipc; // @[Decode.scala 200:27]
  wire [5:0] inst_type = {type_r,type_i,type_s,type_b,type_u,jal}; // @[Cat.scala 30:58]
  wire [51:0] imm_i_hi = io_inst[31] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 72:12]
  wire [11:0] imm_i_lo = io_inst[31:20]; // @[Decode.scala 206:45]
  wire [63:0] imm_i = {imm_i_hi,imm_i_lo}; // @[Cat.scala 30:58]
  wire [6:0] imm_s_hi_lo = io_inst[31:25]; // @[Decode.scala 207:45]
  wire [4:0] imm_s_lo = io_inst[11:7]; // @[Decode.scala 207:59]
  wire [63:0] imm_s = {imm_i_hi,imm_s_hi_lo,imm_s_lo}; // @[Cat.scala 30:58]
  wire [50:0] imm_b_hi_hi_hi = io_inst[31] ? 51'h7ffffffffffff : 51'h0; // @[Bitwise.scala 72:12]
  wire  imm_b_hi_lo = io_inst[7]; // @[Decode.scala 208:55]
  wire [5:0] imm_b_lo_hi_hi = io_inst[30:25]; // @[Decode.scala 208:64]
  wire [3:0] imm_b_lo_hi_lo = io_inst[11:8]; // @[Decode.scala 208:78]
  wire [63:0] imm_b = {imm_b_hi_hi_hi,io_inst[31],imm_b_hi_lo,imm_b_lo_hi_hi,imm_b_lo_hi_lo,1'h0}; // @[Cat.scala 30:58]
  wire [31:0] imm_u_hi_hi = io_inst[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [19:0] imm_u_hi_lo = io_inst[31:12]; // @[Decode.scala 209:45]
  wire [63:0] imm_u = {imm_u_hi_hi,imm_u_hi_lo,12'h0}; // @[Cat.scala 30:58]
  wire [42:0] imm_j_hi_hi_hi = io_inst[31] ? 43'h7ffffffffff : 43'h0; // @[Bitwise.scala 72:12]
  wire [7:0] imm_j_hi_lo = io_inst[19:12]; // @[Decode.scala 210:55]
  wire  imm_j_lo_hi_hi = io_inst[20]; // @[Decode.scala 210:69]
  wire [9:0] imm_j_lo_hi_lo = io_inst[30:21]; // @[Decode.scala 210:79]
  wire [63:0] imm_j = {imm_j_hi_hi_hi,io_inst[31],imm_j_hi_lo,imm_j_lo_hi_hi,imm_j_lo_hi_lo,1'h0}; // @[Cat.scala 30:58]
  wire [63:0] _imm_T_3 = 6'h10 == inst_type ? imm_i : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _imm_T_5 = 6'h8 == inst_type ? imm_s : _imm_T_3; // @[Mux.scala 80:57]
  wire [63:0] _imm_T_7 = 6'h4 == inst_type ? imm_b : _imm_T_5; // @[Mux.scala 80:57]
  wire [63:0] _imm_T_9 = 6'h2 == inst_type ? imm_u : _imm_T_7; // @[Mux.scala 80:57]
  wire [63:0] imm = 6'h1 == inst_type ? imm_j : _imm_T_9; // @[Mux.scala 80:57]
  wire  _io_rs1_en_T = type_r | type_i; // @[Decode.scala 234:25]
  wire [63:0] _bu_jump_pc_T_2 = io_op1 + io_op2; // @[Decode.scala 246:59]
  wire [63:0] _bu_jump_pc_T_3 = _bu_jump_pc_T_2 & 64'hfffffffffffffffe; // @[Decode.scala 246:66]
  wire [63:0] _bu_jump_pc_T_5 = io_pc + imm; // @[Decode.scala 246:95]
  wire [63:0] bu_jump_pc = bu_code == 8'h80 ? _bu_jump_pc_T_3 : _bu_jump_pc_T_5; // @[Decode.scala 246:25]
  wire  _bu_jump_en_T = io_op1 == io_op2; // @[Decode.scala 248:31]
  wire  _bu_jump_en_T_1 = io_op1 != io_op2; // @[Decode.scala 249:31]
  wire  _bu_jump_en_T_4 = $signed(io_op1) < $signed(io_op2); // @[Decode.scala 250:41]
  wire  _bu_jump_en_T_7 = $signed(io_op1) >= $signed(io_op2); // @[Decode.scala 251:41]
  wire  _bu_jump_en_T_8 = io_op1 < io_op2; // @[Decode.scala 252:32]
  wire  _bu_jump_en_T_9 = io_op1 >= io_op2; // @[Decode.scala 253:32]
  wire  _bu_jump_en_T_13 = 8'h2 == bu_code ? _bu_jump_en_T_1 : 8'h1 == bu_code & _bu_jump_en_T; // @[Mux.scala 80:57]
  wire  _bu_jump_en_T_15 = 8'h4 == bu_code ? _bu_jump_en_T_4 : _bu_jump_en_T_13; // @[Mux.scala 80:57]
  wire  _bu_jump_en_T_17 = 8'h8 == bu_code ? _bu_jump_en_T_7 : _bu_jump_en_T_15; // @[Mux.scala 80:57]
  wire  _bu_jump_en_T_19 = 8'h10 == bu_code ? _bu_jump_en_T_8 : _bu_jump_en_T_17; // @[Mux.scala 80:57]
  wire  _bu_jump_en_T_21 = 8'h20 == bu_code ? _bu_jump_en_T_9 : _bu_jump_en_T_19; // @[Mux.scala 80:57]
  wire  bu_jump_en = 8'h80 == bu_code | (8'h40 == bu_code | _bu_jump_en_T_21); // @[Mux.scala 80:57]
  wire [63:0] _csru_jump_pc_T_1 = 8'h1 == csru_code ? io_mtvec : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] csru_jump_pc = 8'h2 == csru_code ? io_mepc : _csru_jump_pc_T_1; // @[Mux.scala 80:57]
  wire  csru_jump_en = 8'h2 == csru_code | 8'h1 == csru_code; // @[Mux.scala 80:57]
  assign io_rs1_en = type_r | type_i | type_s | type_b; // @[Decode.scala 234:45]
  assign io_rs2_en = type_r | type_s | type_b; // @[Decode.scala 235:35]
  assign io_rs1_addr = io_inst[19:15]; // @[Decode.scala 230:24]
  assign io_rs2_addr = io_inst[24:20]; // @[Decode.scala 231:24]
  assign io_rd_en = _io_rs1_en_T | type_u | jal; // @[Decode.scala 236:45]
  assign io_rd_addr = io_inst[11:7]; // @[Decode.scala 232:24]
  assign io_decode_info_fu_code = {fu_code_hi,fu_code_lo}; // @[Cat.scala 30:58]
  assign io_decode_info_alu_code = {alu_code_hi,alu_code_lo}; // @[Cat.scala 30:58]
  assign io_decode_info_bu_code = {bu_code_hi,bu_code_lo}; // @[Cat.scala 30:58]
  assign io_decode_info_lu_code = {lu_code_hi,lu_code_lo}; // @[Cat.scala 30:58]
  assign io_decode_info_su_code = {su_code_hi,su_code_lo}; // @[Cat.scala 30:58]
  assign io_decode_info_mu_code = {mulw,mul}; // @[Cat.scala 30:58]
  assign io_decode_info_du_code = {du_code_hi,du_code_lo}; // @[Cat.scala 30:58]
  assign io_decode_info_csru_code = {csru_code_hi,csru_code_lo}; // @[Cat.scala 30:58]
  assign io_jump_en = bu_jump_en | csru_jump_en; // @[Decode.scala 267:30]
  assign io_jump_pc = bu_jump_en ? bu_jump_pc : csru_jump_pc; // @[Decode.scala 268:22]
  assign io_op1 = io_rs1_en ? io_rs1_data : 64'h0; // @[Decode.scala 238:18]
  assign io_op2 = io_rs2_en ? io_rs2_data : imm; // @[Decode.scala 239:18]
  assign io_imm = 6'h1 == inst_type ? imm_j : _imm_T_9; // @[Mux.scala 80:57]
  assign io_putch = io_inst == 32'h7b; // @[Decode.scala 134:24]
endmodule
module Execution(
  input  [15:0] io_alu_code,
  input  [7:0]  io_bu_code,
  input  [7:0]  io_du_code,
  input  [7:0]  io_csru_code,
  input  [63:0] io_op1,
  input  [63:0] io_op2,
  input  [63:0] io_pc,
  output [63:0] io_alu_out,
  output [63:0] io_bu_out,
  output [63:0] io_du_out,
  output [63:0] io_csru_out,
  input  [4:0]  io_rs1_addr,
  output [11:0] io_csr_raddr,
  input  [63:0] io_csr_rdata,
  output        io_csr_wen,
  output [11:0] io_csr_waddr,
  output [63:0] io_csr_wdata
);
  wire [63:0] _alu_out_T_1 = io_op1 + io_op2; // @[Execution.scala 58:39]
  wire [31:0] alu_out_hi = _alu_out_T_1[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] alu_out_lo = _alu_out_T_1[31:0]; // @[Execution.scala 48:41]
  wire [63:0] _alu_out_T_6 = {alu_out_hi,alu_out_lo}; // @[Cat.scala 30:58]
  wire [63:0] _alu_out_T_8 = io_op1 - io_op2; // @[Execution.scala 60:39]
  wire [31:0] alu_out_hi_1 = _alu_out_T_8[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] alu_out_lo_1 = _alu_out_T_8[31:0]; // @[Execution.scala 48:41]
  wire [63:0] _alu_out_T_13 = {alu_out_hi_1,alu_out_lo_1}; // @[Cat.scala 30:58]
  wire [63:0] _alu_out_T_15 = io_op2 + io_pc; // @[Execution.scala 62:39]
  wire [126:0] _GEN_0 = {{63'd0}, io_op1}; // @[Execution.scala 63:39]
  wire [126:0] _alu_out_T_17 = _GEN_0 << io_op2[5:0]; // @[Execution.scala 63:39]
  wire [63:0] _alu_out_T_20 = io_op1 >> io_op2[5:0]; // @[Execution.scala 64:39]
  wire [63:0] _alu_out_T_24 = $signed(io_op1) >>> io_op2[5:0]; // @[Execution.scala 65:68]
  wire [62:0] _GEN_1 = {{31'd0}, io_op1[31:0]}; // @[Execution.scala 66:51]
  wire [62:0] _alu_out_T_27 = _GEN_1 << io_op2[4:0]; // @[Execution.scala 66:51]
  wire [31:0] alu_out_hi_2 = _alu_out_T_27[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] alu_out_lo_2 = _alu_out_T_27[31:0]; // @[Execution.scala 48:41]
  wire [63:0] _alu_out_T_30 = {alu_out_hi_2,alu_out_lo_2}; // @[Cat.scala 30:58]
  wire [31:0] alu_out_lo_3 = io_op1[31:0] >> io_op2[4:0]; // @[Execution.scala 67:51]
  wire [31:0] alu_out_hi_3 = alu_out_lo_3[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _alu_out_T_36 = {alu_out_hi_3,alu_out_lo_3}; // @[Cat.scala 30:58]
  wire [31:0] _alu_out_T_38 = io_op1[31:0]; // @[Execution.scala 68:57]
  wire [31:0] alu_out_lo_4 = $signed(_alu_out_T_38) >>> io_op2[4:0]; // @[Execution.scala 68:80]
  wire [31:0] alu_out_hi_4 = alu_out_lo_4[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _alu_out_T_44 = {alu_out_hi_4,alu_out_lo_4}; // @[Cat.scala 30:58]
  wire [63:0] _alu_out_T_45 = io_op1 ^ io_op2; // @[Execution.scala 69:39]
  wire [63:0] _alu_out_T_46 = io_op1 | io_op2; // @[Execution.scala 70:39]
  wire [63:0] _alu_out_T_47 = io_op1 & io_op2; // @[Execution.scala 71:39]
  wire  _alu_out_T_50 = $signed(io_op1) < $signed(io_op2); // @[Execution.scala 72:48]
  wire  _alu_out_T_51 = io_op1 < io_op2; // @[Execution.scala 73:39]
  wire [63:0] _alu_out_T_53 = 16'h1 == io_alu_code ? _alu_out_T_1 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _alu_out_T_55 = 16'h2 == io_alu_code ? _alu_out_T_6 : _alu_out_T_53; // @[Mux.scala 80:57]
  wire [63:0] _alu_out_T_57 = 16'h4 == io_alu_code ? _alu_out_T_8 : _alu_out_T_55; // @[Mux.scala 80:57]
  wire [63:0] _alu_out_T_59 = 16'h8 == io_alu_code ? _alu_out_T_13 : _alu_out_T_57; // @[Mux.scala 80:57]
  wire [63:0] _alu_out_T_61 = 16'h10 == io_alu_code ? _alu_out_T_15 : _alu_out_T_59; // @[Mux.scala 80:57]
  wire [63:0] _alu_out_T_63 = 16'h20 == io_alu_code ? _alu_out_T_17[63:0] : _alu_out_T_61; // @[Mux.scala 80:57]
  wire [63:0] _alu_out_T_65 = 16'h40 == io_alu_code ? _alu_out_T_20 : _alu_out_T_63; // @[Mux.scala 80:57]
  wire [63:0] _alu_out_T_67 = 16'h80 == io_alu_code ? _alu_out_T_24 : _alu_out_T_65; // @[Mux.scala 80:57]
  wire [63:0] _alu_out_T_69 = 16'h100 == io_alu_code ? _alu_out_T_30 : _alu_out_T_67; // @[Mux.scala 80:57]
  wire [63:0] _alu_out_T_71 = 16'h200 == io_alu_code ? _alu_out_T_36 : _alu_out_T_69; // @[Mux.scala 80:57]
  wire [63:0] _alu_out_T_73 = 16'h400 == io_alu_code ? _alu_out_T_44 : _alu_out_T_71; // @[Mux.scala 80:57]
  wire [63:0] _alu_out_T_75 = 16'h800 == io_alu_code ? _alu_out_T_45 : _alu_out_T_73; // @[Mux.scala 80:57]
  wire [63:0] _alu_out_T_77 = 16'h1000 == io_alu_code ? _alu_out_T_46 : _alu_out_T_75; // @[Mux.scala 80:57]
  wire [63:0] _alu_out_T_79 = 16'h2000 == io_alu_code ? _alu_out_T_47 : _alu_out_T_77; // @[Mux.scala 80:57]
  wire [63:0] _alu_out_T_81 = 16'h4000 == io_alu_code ? {{63'd0}, _alu_out_T_50} : _alu_out_T_79; // @[Mux.scala 80:57]
  wire [63:0] _bu_out_T_4 = io_pc + 64'h4; // @[Execution.scala 77:81]
  wire [64:0] _du_out_T_3 = $signed(io_op1) / $signed(io_op2); // @[Execution.scala 81:62]
  wire [31:0] _du_out_T_7 = io_op2[31:0]; // @[Execution.scala 82:66]
  wire [32:0] _du_out_T_9 = $signed(_alu_out_T_38) / $signed(_du_out_T_7); // @[Execution.scala 82:76]
  wire [63:0] _du_out_T_10 = io_op1 / io_op2; // @[Execution.scala 83:31]
  wire [31:0] _du_out_T_13 = io_op1[31:0] / io_op2[31:0]; // @[Execution.scala 84:38]
  wire [63:0] _du_out_T_17 = $signed(io_op1) % $signed(io_op2); // @[Execution.scala 85:62]
  wire [31:0] _du_out_T_23 = $signed(_alu_out_T_38) % $signed(_du_out_T_7); // @[Execution.scala 86:76]
  wire [63:0] _GEN_2 = io_op1 % io_op2; // @[Execution.scala 87:31]
  wire [63:0] _du_out_T_24 = _GEN_2[63:0]; // @[Execution.scala 87:31]
  wire [31:0] _GEN_3 = io_op1[31:0] % io_op2[31:0]; // @[Execution.scala 88:38]
  wire [31:0] _du_out_T_27 = _GEN_3[31:0]; // @[Execution.scala 88:38]
  wire [64:0] _du_out_T_29 = 8'h1 == io_du_code ? _du_out_T_3 : 65'h0; // @[Mux.scala 80:57]
  wire [64:0] _du_out_T_31 = 8'h2 == io_du_code ? {{32'd0}, _du_out_T_9} : _du_out_T_29; // @[Mux.scala 80:57]
  wire [64:0] _du_out_T_33 = 8'h4 == io_du_code ? {{1'd0}, _du_out_T_10} : _du_out_T_31; // @[Mux.scala 80:57]
  wire [64:0] _du_out_T_35 = 8'h8 == io_du_code ? {{33'd0}, _du_out_T_13} : _du_out_T_33; // @[Mux.scala 80:57]
  wire [64:0] _du_out_T_37 = 8'h10 == io_du_code ? {{1'd0}, _du_out_T_17} : _du_out_T_35; // @[Mux.scala 80:57]
  wire [64:0] _du_out_T_39 = 8'h20 == io_du_code ? {{33'd0}, _du_out_T_23} : _du_out_T_37; // @[Mux.scala 80:57]
  wire [64:0] _du_out_T_41 = 8'h40 == io_du_code ? {{1'd0}, _du_out_T_24} : _du_out_T_39; // @[Mux.scala 80:57]
  wire [64:0] du_out = 8'h80 == io_du_code ? {{33'd0}, _du_out_T_27} : _du_out_T_41; // @[Mux.scala 80:57]
  wire [63:0] _csru_out_T_1 = 8'h4 == io_csru_code ? io_csr_rdata : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _csru_out_T_3 = 8'h8 == io_csru_code ? io_csr_rdata : _csru_out_T_1; // @[Mux.scala 80:57]
  wire [63:0] _csru_out_T_5 = 8'h10 == io_csru_code ? io_csr_rdata : _csru_out_T_3; // @[Mux.scala 80:57]
  wire [63:0] _csru_out_T_7 = 8'h20 == io_csru_code ? io_csr_rdata : _csru_out_T_5; // @[Mux.scala 80:57]
  wire [63:0] _csru_out_T_9 = 8'h40 == io_csru_code ? io_csr_rdata : _csru_out_T_7; // @[Mux.scala 80:57]
  wire [63:0] _csr_waddr_T_1 = 8'h4 == io_csru_code ? io_op2 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _csr_waddr_T_3 = 8'h8 == io_csru_code ? io_op2 : _csr_waddr_T_1; // @[Mux.scala 80:57]
  wire [63:0] _csr_waddr_T_5 = 8'h10 == io_csru_code ? io_op2 : _csr_waddr_T_3; // @[Mux.scala 80:57]
  wire [63:0] _csr_waddr_T_7 = 8'h20 == io_csru_code ? io_op2 : _csr_waddr_T_5; // @[Mux.scala 80:57]
  wire [63:0] _csr_waddr_T_9 = 8'h40 == io_csru_code ? io_op2 : _csr_waddr_T_7; // @[Mux.scala 80:57]
  wire [63:0] csr_waddr = 8'h80 == io_csru_code ? io_op2 : _csr_waddr_T_9; // @[Mux.scala 80:57]
  wire [63:0] _csr_wdata_T = io_csr_rdata | io_op1; // @[Execution.scala 118:40]
  wire [63:0] _csr_wdata_T_1 = ~io_op1; // @[Execution.scala 120:43]
  wire [63:0] _csr_wdata_T_2 = io_csr_rdata & _csr_wdata_T_1; // @[Execution.scala 120:40]
  wire [63:0] _csr_wdata_T_3 = {59'h0,io_rs1_addr}; // @[Cat.scala 30:58]
  wire [63:0] _csr_wdata_T_4 = io_csr_rdata | _csr_wdata_T_3; // @[Execution.scala 121:40]
  wire [63:0] _csr_wdata_T_7 = ~_csr_wdata_T_3; // @[Execution.scala 123:43]
  wire [63:0] _csr_wdata_T_8 = io_csr_rdata & _csr_wdata_T_7; // @[Execution.scala 123:40]
  wire [63:0] _csr_wdata_T_10 = 8'h4 == io_csru_code ? _csr_wdata_T : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _csr_wdata_T_12 = 8'h8 == io_csru_code ? io_op1 : _csr_wdata_T_10; // @[Mux.scala 80:57]
  wire [63:0] _csr_wdata_T_14 = 8'h10 == io_csru_code ? _csr_wdata_T_2 : _csr_wdata_T_12; // @[Mux.scala 80:57]
  wire [63:0] _csr_wdata_T_16 = 8'h20 == io_csru_code ? _csr_wdata_T_4 : _csr_wdata_T_14; // @[Mux.scala 80:57]
  wire [63:0] _csr_wdata_T_18 = 8'h40 == io_csru_code ? _csr_wdata_T_3 : _csr_wdata_T_16; // @[Mux.scala 80:57]
  assign io_alu_out = 16'h8000 == io_alu_code ? {{63'd0}, _alu_out_T_51} : _alu_out_T_81; // @[Mux.scala 80:57]
  assign io_bu_out = io_bu_code == 8'h80 | io_bu_code == 8'h40 ? _bu_out_T_4 : 64'h0; // @[Execution.scala 77:21]
  assign io_du_out = du_out[63:0]; // @[Execution.scala 129:17]
  assign io_csru_out = 8'h80 == io_csru_code ? io_csr_rdata : _csru_out_T_9; // @[Mux.scala 80:57]
  assign io_csr_raddr = io_op2[11:0]; // @[Execution.scala 92:18]
  assign io_csr_wen = 8'h80 == io_csru_code | (8'h40 == io_csru_code | (8'h20 == io_csru_code | (8'h10 == io_csru_code
     | (8'h8 == io_csru_code | 8'h4 == io_csru_code)))); // @[Mux.scala 80:57]
  assign io_csr_waddr = csr_waddr[11:0]; // @[Execution.scala 134:21]
  assign io_csr_wdata = 8'h80 == io_csru_code ? _csr_wdata_T_8 : _csr_wdata_T_18; // @[Mux.scala 80:57]
endmodule
module RegFile(
  input         clock,
  input         reset,
  input  [4:0]  io_rs1_addr,
  input  [4:0]  io_rs2_addr,
  output [63:0] io_rs1_data,
  output [63:0] io_rs2_data,
  input  [4:0]  io_rd_addr,
  input  [63:0] io_rd_data,
  input         io_rd_en,
  output [63:0] rf_10
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  wire  dt_ar_clock; // @[RegFile.scala 27:23]
  wire [7:0] dt_ar_coreid; // @[RegFile.scala 27:23]
  wire [63:0] dt_ar_gpr_0; // @[RegFile.scala 27:23]
  wire [63:0] dt_ar_gpr_1; // @[RegFile.scala 27:23]
  wire [63:0] dt_ar_gpr_2; // @[RegFile.scala 27:23]
  wire [63:0] dt_ar_gpr_3; // @[RegFile.scala 27:23]
  wire [63:0] dt_ar_gpr_4; // @[RegFile.scala 27:23]
  wire [63:0] dt_ar_gpr_5; // @[RegFile.scala 27:23]
  wire [63:0] dt_ar_gpr_6; // @[RegFile.scala 27:23]
  wire [63:0] dt_ar_gpr_7; // @[RegFile.scala 27:23]
  wire [63:0] dt_ar_gpr_8; // @[RegFile.scala 27:23]
  wire [63:0] dt_ar_gpr_9; // @[RegFile.scala 27:23]
  wire [63:0] dt_ar_gpr_10; // @[RegFile.scala 27:23]
  wire [63:0] dt_ar_gpr_11; // @[RegFile.scala 27:23]
  wire [63:0] dt_ar_gpr_12; // @[RegFile.scala 27:23]
  wire [63:0] dt_ar_gpr_13; // @[RegFile.scala 27:23]
  wire [63:0] dt_ar_gpr_14; // @[RegFile.scala 27:23]
  wire [63:0] dt_ar_gpr_15; // @[RegFile.scala 27:23]
  wire [63:0] dt_ar_gpr_16; // @[RegFile.scala 27:23]
  wire [63:0] dt_ar_gpr_17; // @[RegFile.scala 27:23]
  wire [63:0] dt_ar_gpr_18; // @[RegFile.scala 27:23]
  wire [63:0] dt_ar_gpr_19; // @[RegFile.scala 27:23]
  wire [63:0] dt_ar_gpr_20; // @[RegFile.scala 27:23]
  wire [63:0] dt_ar_gpr_21; // @[RegFile.scala 27:23]
  wire [63:0] dt_ar_gpr_22; // @[RegFile.scala 27:23]
  wire [63:0] dt_ar_gpr_23; // @[RegFile.scala 27:23]
  wire [63:0] dt_ar_gpr_24; // @[RegFile.scala 27:23]
  wire [63:0] dt_ar_gpr_25; // @[RegFile.scala 27:23]
  wire [63:0] dt_ar_gpr_26; // @[RegFile.scala 27:23]
  wire [63:0] dt_ar_gpr_27; // @[RegFile.scala 27:23]
  wire [63:0] dt_ar_gpr_28; // @[RegFile.scala 27:23]
  wire [63:0] dt_ar_gpr_29; // @[RegFile.scala 27:23]
  wire [63:0] dt_ar_gpr_30; // @[RegFile.scala 27:23]
  wire [63:0] dt_ar_gpr_31; // @[RegFile.scala 27:23]
  reg [63:0] rf__0; // @[RegFile.scala 16:19]
  reg [63:0] rf__1; // @[RegFile.scala 16:19]
  reg [63:0] rf__2; // @[RegFile.scala 16:19]
  reg [63:0] rf__3; // @[RegFile.scala 16:19]
  reg [63:0] rf__4; // @[RegFile.scala 16:19]
  reg [63:0] rf__5; // @[RegFile.scala 16:19]
  reg [63:0] rf__6; // @[RegFile.scala 16:19]
  reg [63:0] rf__7; // @[RegFile.scala 16:19]
  reg [63:0] rf__8; // @[RegFile.scala 16:19]
  reg [63:0] rf__9; // @[RegFile.scala 16:19]
  reg [63:0] rf__10; // @[RegFile.scala 16:19]
  reg [63:0] rf__11; // @[RegFile.scala 16:19]
  reg [63:0] rf__12; // @[RegFile.scala 16:19]
  reg [63:0] rf__13; // @[RegFile.scala 16:19]
  reg [63:0] rf__14; // @[RegFile.scala 16:19]
  reg [63:0] rf__15; // @[RegFile.scala 16:19]
  reg [63:0] rf__16; // @[RegFile.scala 16:19]
  reg [63:0] rf__17; // @[RegFile.scala 16:19]
  reg [63:0] rf__18; // @[RegFile.scala 16:19]
  reg [63:0] rf__19; // @[RegFile.scala 16:19]
  reg [63:0] rf__20; // @[RegFile.scala 16:19]
  reg [63:0] rf__21; // @[RegFile.scala 16:19]
  reg [63:0] rf__22; // @[RegFile.scala 16:19]
  reg [63:0] rf__23; // @[RegFile.scala 16:19]
  reg [63:0] rf__24; // @[RegFile.scala 16:19]
  reg [63:0] rf__25; // @[RegFile.scala 16:19]
  reg [63:0] rf__26; // @[RegFile.scala 16:19]
  reg [63:0] rf__27; // @[RegFile.scala 16:19]
  reg [63:0] rf__28; // @[RegFile.scala 16:19]
  reg [63:0] rf__29; // @[RegFile.scala 16:19]
  reg [63:0] rf__30; // @[RegFile.scala 16:19]
  reg [63:0] rf__31; // @[RegFile.scala 16:19]
  wire [63:0] _GEN_65 = 5'h1 == io_rs1_addr ? rf__1 : rf__0; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_66 = 5'h2 == io_rs1_addr ? rf__2 : _GEN_65; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_67 = 5'h3 == io_rs1_addr ? rf__3 : _GEN_66; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_68 = 5'h4 == io_rs1_addr ? rf__4 : _GEN_67; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_69 = 5'h5 == io_rs1_addr ? rf__5 : _GEN_68; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_70 = 5'h6 == io_rs1_addr ? rf__6 : _GEN_69; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_71 = 5'h7 == io_rs1_addr ? rf__7 : _GEN_70; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_72 = 5'h8 == io_rs1_addr ? rf__8 : _GEN_71; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_73 = 5'h9 == io_rs1_addr ? rf__9 : _GEN_72; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_74 = 5'ha == io_rs1_addr ? rf__10 : _GEN_73; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_75 = 5'hb == io_rs1_addr ? rf__11 : _GEN_74; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_76 = 5'hc == io_rs1_addr ? rf__12 : _GEN_75; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_77 = 5'hd == io_rs1_addr ? rf__13 : _GEN_76; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_78 = 5'he == io_rs1_addr ? rf__14 : _GEN_77; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_79 = 5'hf == io_rs1_addr ? rf__15 : _GEN_78; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_80 = 5'h10 == io_rs1_addr ? rf__16 : _GEN_79; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_81 = 5'h11 == io_rs1_addr ? rf__17 : _GEN_80; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_82 = 5'h12 == io_rs1_addr ? rf__18 : _GEN_81; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_83 = 5'h13 == io_rs1_addr ? rf__19 : _GEN_82; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_84 = 5'h14 == io_rs1_addr ? rf__20 : _GEN_83; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_85 = 5'h15 == io_rs1_addr ? rf__21 : _GEN_84; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_86 = 5'h16 == io_rs1_addr ? rf__22 : _GEN_85; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_87 = 5'h17 == io_rs1_addr ? rf__23 : _GEN_86; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_88 = 5'h18 == io_rs1_addr ? rf__24 : _GEN_87; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_89 = 5'h19 == io_rs1_addr ? rf__25 : _GEN_88; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_90 = 5'h1a == io_rs1_addr ? rf__26 : _GEN_89; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_91 = 5'h1b == io_rs1_addr ? rf__27 : _GEN_90; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_92 = 5'h1c == io_rs1_addr ? rf__28 : _GEN_91; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_93 = 5'h1d == io_rs1_addr ? rf__29 : _GEN_92; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_94 = 5'h1e == io_rs1_addr ? rf__30 : _GEN_93; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_95 = 5'h1f == io_rs1_addr ? rf__31 : _GEN_94; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_97 = 5'h1 == io_rs2_addr ? rf__1 : rf__0; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_98 = 5'h2 == io_rs2_addr ? rf__2 : _GEN_97; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_99 = 5'h3 == io_rs2_addr ? rf__3 : _GEN_98; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_100 = 5'h4 == io_rs2_addr ? rf__4 : _GEN_99; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_101 = 5'h5 == io_rs2_addr ? rf__5 : _GEN_100; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_102 = 5'h6 == io_rs2_addr ? rf__6 : _GEN_101; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_103 = 5'h7 == io_rs2_addr ? rf__7 : _GEN_102; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_104 = 5'h8 == io_rs2_addr ? rf__8 : _GEN_103; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_105 = 5'h9 == io_rs2_addr ? rf__9 : _GEN_104; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_106 = 5'ha == io_rs2_addr ? rf__10 : _GEN_105; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_107 = 5'hb == io_rs2_addr ? rf__11 : _GEN_106; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_108 = 5'hc == io_rs2_addr ? rf__12 : _GEN_107; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_109 = 5'hd == io_rs2_addr ? rf__13 : _GEN_108; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_110 = 5'he == io_rs2_addr ? rf__14 : _GEN_109; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_111 = 5'hf == io_rs2_addr ? rf__15 : _GEN_110; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_112 = 5'h10 == io_rs2_addr ? rf__16 : _GEN_111; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_113 = 5'h11 == io_rs2_addr ? rf__17 : _GEN_112; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_114 = 5'h12 == io_rs2_addr ? rf__18 : _GEN_113; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_115 = 5'h13 == io_rs2_addr ? rf__19 : _GEN_114; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_116 = 5'h14 == io_rs2_addr ? rf__20 : _GEN_115; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_117 = 5'h15 == io_rs2_addr ? rf__21 : _GEN_116; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_118 = 5'h16 == io_rs2_addr ? rf__22 : _GEN_117; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_119 = 5'h17 == io_rs2_addr ? rf__23 : _GEN_118; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_120 = 5'h18 == io_rs2_addr ? rf__24 : _GEN_119; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_121 = 5'h19 == io_rs2_addr ? rf__25 : _GEN_120; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_122 = 5'h1a == io_rs2_addr ? rf__26 : _GEN_121; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_123 = 5'h1b == io_rs2_addr ? rf__27 : _GEN_122; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_124 = 5'h1c == io_rs2_addr ? rf__28 : _GEN_123; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_125 = 5'h1d == io_rs2_addr ? rf__29 : _GEN_124; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_126 = 5'h1e == io_rs2_addr ? rf__30 : _GEN_125; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_127 = 5'h1f == io_rs2_addr ? rf__31 : _GEN_126; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  DifftestArchIntRegState dt_ar ( // @[RegFile.scala 27:23]
    .clock(dt_ar_clock),
    .coreid(dt_ar_coreid),
    .gpr_0(dt_ar_gpr_0),
    .gpr_1(dt_ar_gpr_1),
    .gpr_2(dt_ar_gpr_2),
    .gpr_3(dt_ar_gpr_3),
    .gpr_4(dt_ar_gpr_4),
    .gpr_5(dt_ar_gpr_5),
    .gpr_6(dt_ar_gpr_6),
    .gpr_7(dt_ar_gpr_7),
    .gpr_8(dt_ar_gpr_8),
    .gpr_9(dt_ar_gpr_9),
    .gpr_10(dt_ar_gpr_10),
    .gpr_11(dt_ar_gpr_11),
    .gpr_12(dt_ar_gpr_12),
    .gpr_13(dt_ar_gpr_13),
    .gpr_14(dt_ar_gpr_14),
    .gpr_15(dt_ar_gpr_15),
    .gpr_16(dt_ar_gpr_16),
    .gpr_17(dt_ar_gpr_17),
    .gpr_18(dt_ar_gpr_18),
    .gpr_19(dt_ar_gpr_19),
    .gpr_20(dt_ar_gpr_20),
    .gpr_21(dt_ar_gpr_21),
    .gpr_22(dt_ar_gpr_22),
    .gpr_23(dt_ar_gpr_23),
    .gpr_24(dt_ar_gpr_24),
    .gpr_25(dt_ar_gpr_25),
    .gpr_26(dt_ar_gpr_26),
    .gpr_27(dt_ar_gpr_27),
    .gpr_28(dt_ar_gpr_28),
    .gpr_29(dt_ar_gpr_29),
    .gpr_30(dt_ar_gpr_30),
    .gpr_31(dt_ar_gpr_31)
  );
  assign io_rs1_data = io_rs1_addr != 5'h0 ? _GEN_95 : 64'h0; // @[RegFile.scala 22:21]
  assign io_rs2_data = io_rs2_addr != 5'h0 ? _GEN_127 : 64'h0; // @[RegFile.scala 23:21]
  assign rf_10 = rf__10;
  assign dt_ar_clock = clock; // @[RegFile.scala 28:21]
  assign dt_ar_coreid = 8'h0; // @[RegFile.scala 29:21]
  assign dt_ar_gpr_0 = rf__0; // @[RegFile.scala 30:21]
  assign dt_ar_gpr_1 = rf__1; // @[RegFile.scala 30:21]
  assign dt_ar_gpr_2 = rf__2; // @[RegFile.scala 30:21]
  assign dt_ar_gpr_3 = rf__3; // @[RegFile.scala 30:21]
  assign dt_ar_gpr_4 = rf__4; // @[RegFile.scala 30:21]
  assign dt_ar_gpr_5 = rf__5; // @[RegFile.scala 30:21]
  assign dt_ar_gpr_6 = rf__6; // @[RegFile.scala 30:21]
  assign dt_ar_gpr_7 = rf__7; // @[RegFile.scala 30:21]
  assign dt_ar_gpr_8 = rf__8; // @[RegFile.scala 30:21]
  assign dt_ar_gpr_9 = rf__9; // @[RegFile.scala 30:21]
  assign dt_ar_gpr_10 = rf__10; // @[RegFile.scala 30:21]
  assign dt_ar_gpr_11 = rf__11; // @[RegFile.scala 30:21]
  assign dt_ar_gpr_12 = rf__12; // @[RegFile.scala 30:21]
  assign dt_ar_gpr_13 = rf__13; // @[RegFile.scala 30:21]
  assign dt_ar_gpr_14 = rf__14; // @[RegFile.scala 30:21]
  assign dt_ar_gpr_15 = rf__15; // @[RegFile.scala 30:21]
  assign dt_ar_gpr_16 = rf__16; // @[RegFile.scala 30:21]
  assign dt_ar_gpr_17 = rf__17; // @[RegFile.scala 30:21]
  assign dt_ar_gpr_18 = rf__18; // @[RegFile.scala 30:21]
  assign dt_ar_gpr_19 = rf__19; // @[RegFile.scala 30:21]
  assign dt_ar_gpr_20 = rf__20; // @[RegFile.scala 30:21]
  assign dt_ar_gpr_21 = rf__21; // @[RegFile.scala 30:21]
  assign dt_ar_gpr_22 = rf__22; // @[RegFile.scala 30:21]
  assign dt_ar_gpr_23 = rf__23; // @[RegFile.scala 30:21]
  assign dt_ar_gpr_24 = rf__24; // @[RegFile.scala 30:21]
  assign dt_ar_gpr_25 = rf__25; // @[RegFile.scala 30:21]
  assign dt_ar_gpr_26 = rf__26; // @[RegFile.scala 30:21]
  assign dt_ar_gpr_27 = rf__27; // @[RegFile.scala 30:21]
  assign dt_ar_gpr_28 = rf__28; // @[RegFile.scala 30:21]
  assign dt_ar_gpr_29 = rf__29; // @[RegFile.scala 30:21]
  assign dt_ar_gpr_30 = rf__30; // @[RegFile.scala 30:21]
  assign dt_ar_gpr_31 = rf__31; // @[RegFile.scala 30:21]
  always @(posedge clock) begin
    if (reset) begin // @[RegFile.scala 16:19]
      rf__0 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h0 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__0 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__1 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h1 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__1 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__2 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h2 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__2 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__3 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h3 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__3 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__4 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h4 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__4 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__5 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h5 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__5 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__6 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h6 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__6 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__7 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h7 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__7 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__8 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h8 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__8 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__9 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h9 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__9 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__10 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'ha == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__10 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__11 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'hb == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__11 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__12 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'hc == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__12 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__13 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'hd == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__13 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__14 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'he == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__14 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__15 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'hf == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__15 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__16 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h10 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__16 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__17 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h11 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__17 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__18 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h12 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__18 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__19 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h13 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__19 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__20 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h14 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__20 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__21 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h15 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__21 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__22 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h16 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__22 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__23 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h17 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__23 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__24 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h18 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__24 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__25 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h19 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__25 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__26 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h1a == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__26 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__27 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h1b == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__27 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__28 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h1c == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__28 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__29 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h1d == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__29 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__30 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h1e == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__30 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__31 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h1f == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__31 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  rf__0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  rf__1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  rf__2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  rf__3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  rf__4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  rf__5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  rf__6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  rf__7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  rf__8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  rf__9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  rf__10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  rf__11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  rf__12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  rf__13 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  rf__14 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  rf__15 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  rf__16 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  rf__17 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  rf__18 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  rf__19 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  rf__20 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  rf__21 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  rf__22 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  rf__23 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  rf__24 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  rf__25 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  rf__26 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  rf__27 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  rf__28 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  rf__29 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  rf__30 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  rf__31 = _RAND_31[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Csr(
  input         clock,
  input         reset,
  input  [11:0] io_raddr,
  output [63:0] io_rdata,
  input         io_wen,
  input  [11:0] io_waddr,
  input  [63:0] io_wdata,
  input         io_set_mtip,
  input         io_clear_mtip,
  input         io_exception,
  input  [63:0] io_cause,
  input         io_mret,
  input  [63:0] io_pc,
  output [63:0] io_mtvec,
  output [63:0] io_mepc,
  output        io_time_intr
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  dt_cs_clock; // @[Csr.scala 114:27]
  wire [7:0] dt_cs_coreid; // @[Csr.scala 114:27]
  wire [1:0] dt_cs_priviledgeMode; // @[Csr.scala 114:27]
  wire [63:0] dt_cs_mstatus; // @[Csr.scala 114:27]
  wire [63:0] dt_cs_sstatus; // @[Csr.scala 114:27]
  wire [63:0] dt_cs_mepc; // @[Csr.scala 114:27]
  wire [63:0] dt_cs_sepc; // @[Csr.scala 114:27]
  wire [63:0] dt_cs_mtval; // @[Csr.scala 114:27]
  wire [63:0] dt_cs_stval; // @[Csr.scala 114:27]
  wire [63:0] dt_cs_mtvec; // @[Csr.scala 114:27]
  wire [63:0] dt_cs_stvec; // @[Csr.scala 114:27]
  wire [63:0] dt_cs_mcause; // @[Csr.scala 114:27]
  wire [63:0] dt_cs_scause; // @[Csr.scala 114:27]
  wire [63:0] dt_cs_satp; // @[Csr.scala 114:27]
  wire [63:0] dt_cs_mip; // @[Csr.scala 114:27]
  wire [63:0] dt_cs_mie; // @[Csr.scala 114:27]
  wire [63:0] dt_cs_mscratch; // @[Csr.scala 114:27]
  wire [63:0] dt_cs_sscratch; // @[Csr.scala 114:27]
  wire [63:0] dt_cs_mideleg; // @[Csr.scala 114:27]
  wire [63:0] dt_cs_medeleg; // @[Csr.scala 114:27]
  reg [63:0] mstatus; // @[Csr.scala 44:30]
  reg [63:0] mtvec; // @[Csr.scala 45:30]
  reg [63:0] mepc; // @[Csr.scala 46:30]
  reg [63:0] mcause; // @[Csr.scala 47:30]
  reg [63:0] mcycle; // @[Csr.scala 48:30]
  reg [63:0] mhartid; // @[Csr.scala 50:30]
  reg [63:0] mie; // @[Csr.scala 51:30]
  reg [63:0] mip; // @[Csr.scala 52:30]
  reg [63:0] mscratch; // @[Csr.scala 53:30]
  reg [63:0] satp; // @[Csr.scala 54:30]
  wire [63:0] _io_rdata_T_1 = 12'h300 == io_raddr ? mstatus : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _io_rdata_T_3 = 12'h305 == io_raddr ? mtvec : _io_rdata_T_1; // @[Mux.scala 80:57]
  wire [63:0] _io_rdata_T_5 = 12'h341 == io_raddr ? mepc : _io_rdata_T_3; // @[Mux.scala 80:57]
  wire [63:0] _io_rdata_T_7 = 12'h342 == io_raddr ? mcause : _io_rdata_T_5; // @[Mux.scala 80:57]
  wire [63:0] _io_rdata_T_9 = 12'hb00 == io_raddr ? mcycle : _io_rdata_T_7; // @[Mux.scala 80:57]
  wire [63:0] _io_rdata_T_11 = 12'hf14 == io_raddr ? mhartid : _io_rdata_T_9; // @[Mux.scala 80:57]
  wire [63:0] _io_rdata_T_13 = 12'h304 == io_raddr ? mie : _io_rdata_T_11; // @[Mux.scala 80:57]
  wire [63:0] _io_rdata_T_15 = 12'h344 == io_raddr ? mip : _io_rdata_T_13; // @[Mux.scala 80:57]
  wire [63:0] _io_rdata_T_17 = 12'h340 == io_raddr ? mscratch : _io_rdata_T_15; // @[Mux.scala 80:57]
  wire [63:0] _mcycle_T_3 = mcycle + 64'h1; // @[Csr.scala 69:68]
  wire  mstatus_SD = io_wdata[14:13] == 2'h3 | io_wdata[16:15] == 2'h3; // @[Csr.scala 71:60]
  wire [50:0] mstatus_hi_hi_hi = mstatus[63:13]; // @[Csr.scala 74:31]
  wire [2:0] mstatus_hi_lo_hi = mstatus[10:8]; // @[Csr.scala 74:61]
  wire  mstatus_hi_lo_lo = mstatus[3]; // @[Csr.scala 74:76]
  wire [2:0] mstatus_lo_hi_hi = mstatus[6:4]; // @[Csr.scala 74:88]
  wire [2:0] mstatus_lo_lo = mstatus[2:0]; // @[Csr.scala 74:108]
  wire [63:0] _mstatus_T = {mstatus_hi_hi_hi,2'h3,mstatus_hi_lo_hi,mstatus_hi_lo_lo,mstatus_lo_hi_hi,1'h0,mstatus_lo_lo}
    ; // @[Cat.scala 30:58]
  wire  mstatus_lo_hi_lo = mstatus[7]; // @[Csr.scala 77:96]
  wire [63:0] _mstatus_T_1 = {mstatus_hi_hi_hi,2'h0,mstatus_hi_lo_hi,1'h1,mstatus_lo_hi_hi,mstatus_lo_hi_lo,
    mstatus_lo_lo}; // @[Cat.scala 30:58]
  wire [62:0] mstatus_lo_2 = io_wdata[62:0]; // @[Csr.scala 80:44]
  wire [63:0] _mstatus_T_2 = {mstatus_SD,mstatus_lo_2}; // @[Cat.scala 30:58]
  wire [61:0] mepc_hi = io_wdata[63:2]; // @[Csr.scala 89:65]
  wire [63:0] _mepc_T = {mepc_hi,2'h0}; // @[Cat.scala 30:58]
  wire [63:0] _mip_T = mip & 64'hffffffffffffff7f; // @[Csr.scala 96:37]
  wire [63:0] _mip_T_1 = mip | 64'h80; // @[Csr.scala 97:40]
  wire [55:0] mip_hi_hi = io_wdata[63:8]; // @[Csr.scala 98:63]
  wire  mip_hi_lo = mip[7]; // @[Csr.scala 98:75]
  wire [6:0] mip_lo = io_wdata[6:0]; // @[Csr.scala 98:88]
  wire [63:0] _mip_T_2 = {mip_hi_hi,mip_hi_lo,mip_lo}; // @[Cat.scala 30:58]
  DifftestCSRState dt_cs ( // @[Csr.scala 114:27]
    .clock(dt_cs_clock),
    .coreid(dt_cs_coreid),
    .priviledgeMode(dt_cs_priviledgeMode),
    .mstatus(dt_cs_mstatus),
    .sstatus(dt_cs_sstatus),
    .mepc(dt_cs_mepc),
    .sepc(dt_cs_sepc),
    .mtval(dt_cs_mtval),
    .stval(dt_cs_stval),
    .mtvec(dt_cs_mtvec),
    .stvec(dt_cs_stvec),
    .mcause(dt_cs_mcause),
    .scause(dt_cs_scause),
    .satp(dt_cs_satp),
    .mip(dt_cs_mip),
    .mie(dt_cs_mie),
    .mscratch(dt_cs_mscratch),
    .sscratch(dt_cs_sscratch),
    .mideleg(dt_cs_mideleg),
    .medeleg(dt_cs_medeleg)
  );
  assign io_rdata = 12'h180 == io_raddr ? satp : _io_rdata_T_17; // @[Mux.scala 80:57]
  assign io_mtvec = mtvec; // @[Csr.scala 108:14]
  assign io_mepc = mepc; // @[Csr.scala 109:14]
  assign io_time_intr = mip_hi_lo & mie[7] & mstatus_hi_lo_lo; // @[Csr.scala 110:38]
  assign dt_cs_clock = clock; // @[Csr.scala 115:33]
  assign dt_cs_coreid = 8'h0; // @[Csr.scala 116:33]
  assign dt_cs_priviledgeMode = 2'h3; // @[Csr.scala 117:33]
  assign dt_cs_mstatus = mstatus; // @[Csr.scala 118:33]
  assign dt_cs_sstatus = mstatus & 64'h80000003000de122; // @[Csr.scala 119:44]
  assign dt_cs_mepc = mepc; // @[Csr.scala 120:33]
  assign dt_cs_sepc = 64'h0; // @[Csr.scala 121:33]
  assign dt_cs_mtval = 64'h0; // @[Csr.scala 122:33]
  assign dt_cs_stval = 64'h0; // @[Csr.scala 123:33]
  assign dt_cs_mtvec = mtvec; // @[Csr.scala 124:33]
  assign dt_cs_stvec = 64'h0; // @[Csr.scala 125:33]
  assign dt_cs_mcause = mcause; // @[Csr.scala 126:33]
  assign dt_cs_scause = 64'h0; // @[Csr.scala 127:33]
  assign dt_cs_satp = satp; // @[Csr.scala 128:33]
  assign dt_cs_mip = 64'h0;
  assign dt_cs_mie = mie; // @[Csr.scala 130:33]
  assign dt_cs_mscratch = mscratch; // @[Csr.scala 131:33]
  assign dt_cs_sscratch = 64'h0; // @[Csr.scala 132:33]
  assign dt_cs_mideleg = 64'h0; // @[Csr.scala 133:33]
  assign dt_cs_medeleg = 64'h0; // @[Csr.scala 134:33]
  always @(posedge clock) begin
    if (reset) begin // @[Csr.scala 44:30]
      mstatus <= 64'h1800; // @[Csr.scala 44:30]
    end else if (io_exception) begin // @[Csr.scala 73:23]
      mstatus <= _mstatus_T; // @[Csr.scala 74:17]
    end else if (io_mret) begin // @[Csr.scala 76:23]
      mstatus <= _mstatus_T_1; // @[Csr.scala 77:17]
    end else if (io_wen & io_waddr == 12'h300) begin // @[Csr.scala 79:46]
      mstatus <= _mstatus_T_2; // @[Csr.scala 80:17]
    end
    if (reset) begin // @[Csr.scala 45:30]
      mtvec <= 64'h0; // @[Csr.scala 45:30]
    end else if (io_wen & io_waddr == 12'h305) begin // @[Csr.scala 86:17]
      mtvec <= io_wdata;
    end
    if (reset) begin // @[Csr.scala 46:30]
      mepc <= 64'h0; // @[Csr.scala 46:30]
    end else if (io_exception) begin // @[Csr.scala 88:24]
      mepc <= io_pc; // @[Csr.scala 88:30]
    end else if (io_wen & io_waddr == 12'h341) begin // @[Csr.scala 89:44]
      mepc <= _mepc_T; // @[Csr.scala 89:50]
    end
    if (reset) begin // @[Csr.scala 47:30]
      mcause <= 64'h0; // @[Csr.scala 47:30]
    end else if (io_exception) begin // @[Csr.scala 92:24]
      mcause <= io_cause; // @[Csr.scala 92:32]
    end else if (io_wen & io_waddr == 12'h342) begin // @[Csr.scala 93:46]
      mcause <= io_wdata; // @[Csr.scala 93:54]
    end
    if (reset) begin // @[Csr.scala 48:30]
      mcycle <= 64'h0; // @[Csr.scala 48:30]
    end else if (io_wen & io_waddr == 12'hb00) begin // @[Csr.scala 69:19]
      mcycle <= io_wdata;
    end else begin
      mcycle <= _mcycle_T_3;
    end
    if (reset) begin // @[Csr.scala 50:30]
      mhartid <= 64'h0; // @[Csr.scala 50:30]
    end else if (io_wen & io_waddr == 12'hf14) begin // @[Csr.scala 102:23]
      mhartid <= io_wdata;
    end
    if (reset) begin // @[Csr.scala 51:30]
      mie <= 64'h0; // @[Csr.scala 51:30]
    end else if (io_wen & io_waddr == 12'h304) begin // @[Csr.scala 103:23]
      mie <= io_wdata;
    end
    if (reset) begin // @[Csr.scala 52:30]
      mip <= 64'h0; // @[Csr.scala 52:30]
    end else if (io_clear_mtip) begin // @[Csr.scala 96:25]
      mip <= _mip_T; // @[Csr.scala 96:30]
    end else if (io_set_mtip) begin // @[Csr.scala 97:28]
      mip <= _mip_T_1; // @[Csr.scala 97:33]
    end else if (io_wen & io_waddr == 12'h344) begin // @[Csr.scala 98:43]
      mip <= _mip_T_2; // @[Csr.scala 98:48]
    end
    if (reset) begin // @[Csr.scala 53:30]
      mscratch <= 64'h0; // @[Csr.scala 53:30]
    end else if (io_wen & io_waddr == 12'h340) begin // @[Csr.scala 104:23]
      mscratch <= io_wdata;
    end
    if (reset) begin // @[Csr.scala 54:30]
      satp <= 64'h0; // @[Csr.scala 54:30]
    end else if (io_wen & io_waddr == 12'h180) begin // @[Csr.scala 105:23]
      satp <= io_wdata;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mstatus = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  mtvec = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  mepc = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  mcause = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  mcycle = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  mhartid = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  mie = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  mip = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  mscratch = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  satp = _RAND_9[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PreAccessMemory(
  input  [6:0]  io_lu_code,
  input  [3:0]  io_su_code,
  input  [63:0] io_op1,
  input  [63:0] io_op2,
  input  [63:0] io_imm,
  output [5:0]  io_lu_shift,
  output        io_ren,
  output [63:0] io_raddr,
  output        io_wen,
  output [63:0] io_waddr,
  output [63:0] io_wdata,
  output [7:0]  io_wmask,
  output [2:0]  io_transfer
);
  wire [63:0] lu_offset = io_op1 + io_op2; // @[PreAccessMemory.scala 25:28]
  wire [63:0] su_offset = io_op1 + io_imm; // @[PreAccessMemory.scala 31:28]
  wire [5:0] su_shift = {su_offset[2:0], 3'h0}; // @[PreAccessMemory.scala 32:37]
  wire [126:0] _GEN_0 = {{63'd0}, io_op2}; // @[PreAccessMemory.scala 35:28]
  wire [126:0] su_wdata = _GEN_0 << su_shift; // @[PreAccessMemory.scala 35:28]
  wire [7:0] _su_wmask_T_1 = 8'h1 << su_offset[2:0]; // @[PreAccessMemory.scala 37:37]
  wire [8:0] _su_wmask_T_3 = 9'h3 << su_offset[2:0]; // @[PreAccessMemory.scala 38:37]
  wire [10:0] _su_wmask_T_5 = 11'hf << su_offset[2:0]; // @[PreAccessMemory.scala 39:37]
  wire [7:0] _su_wmask_T_7 = 4'h1 == io_su_code ? _su_wmask_T_1 : 8'h0; // @[Mux.scala 80:57]
  wire [8:0] _su_wmask_T_9 = 4'h2 == io_su_code ? _su_wmask_T_3 : {{1'd0}, _su_wmask_T_7}; // @[Mux.scala 80:57]
  wire [10:0] _su_wmask_T_11 = 4'h4 == io_su_code ? _su_wmask_T_5 : {{2'd0}, _su_wmask_T_9}; // @[Mux.scala 80:57]
  wire [10:0] su_wmask = 4'h8 == io_su_code ? 11'hff : _su_wmask_T_11; // @[Mux.scala 80:57]
  wire [10:0] _transfer_T = {io_su_code,io_lu_code}; // @[Cat.scala 30:58]
  wire [1:0] _transfer_T_6 = 11'h4 == _transfer_T ? 2'h2 : {{1'd0}, 11'h2 == _transfer_T}; // @[Mux.scala 80:57]
  wire [1:0] _transfer_T_8 = 11'h8 == _transfer_T ? 2'h3 : _transfer_T_6; // @[Mux.scala 80:57]
  wire [1:0] _transfer_T_10 = 11'h10 == _transfer_T ? 2'h0 : _transfer_T_8; // @[Mux.scala 80:57]
  wire [1:0] _transfer_T_12 = 11'h20 == _transfer_T ? 2'h1 : _transfer_T_10; // @[Mux.scala 80:57]
  wire [1:0] _transfer_T_14 = 11'h40 == _transfer_T ? 2'h2 : _transfer_T_12; // @[Mux.scala 80:57]
  wire [1:0] _transfer_T_16 = 11'h80 == _transfer_T ? 2'h0 : _transfer_T_14; // @[Mux.scala 80:57]
  wire [1:0] _transfer_T_18 = 11'h100 == _transfer_T ? 2'h1 : _transfer_T_16; // @[Mux.scala 80:57]
  wire [1:0] _transfer_T_20 = 11'h200 == _transfer_T ? 2'h2 : _transfer_T_18; // @[Mux.scala 80:57]
  wire [1:0] transfer = 11'h400 == _transfer_T ? 2'h3 : _transfer_T_20; // @[Mux.scala 80:57]
  assign io_lu_shift = {lu_offset[2:0], 3'h0}; // @[PreAccessMemory.scala 26:36]
  assign io_ren = io_lu_code != 7'h0; // @[PreAccessMemory.scala 27:29]
  assign io_raddr = io_op1 + io_op2; // @[PreAccessMemory.scala 25:28]
  assign io_wen = io_su_code != 4'h0; // @[PreAccessMemory.scala 33:32]
  assign io_waddr = io_op1 + io_imm; // @[PreAccessMemory.scala 31:28]
  assign io_wdata = su_wdata[63:0]; // @[PreAccessMemory.scala 63:17]
  assign io_wmask = su_wmask[7:0]; // @[PreAccessMemory.scala 64:17]
  assign io_transfer = {{1'd0}, transfer}; // @[Mux.scala 80:57]
endmodule
module AccessMemory(
  input  [6:0]  io_lu_code,
  input  [5:0]  io_lu_shift,
  input  [63:0] io_rdata,
  output [63:0] io_lu_out
);
  wire [63:0] _io_lu_out_T = io_rdata >> io_lu_shift; // @[AccessMemory.scala 23:41]
  wire [55:0] io_lu_out_hi = _io_lu_out_T[7] ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 72:12]
  wire [7:0] io_lu_out_lo = _io_lu_out_T[7:0]; // @[AccessMemory.scala 13:40]
  wire [63:0] _io_lu_out_T_3 = {io_lu_out_hi,io_lu_out_lo}; // @[Cat.scala 30:58]
  wire [47:0] io_lu_out_hi_1 = _io_lu_out_T[15] ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 72:12]
  wire [15:0] io_lu_out_lo_1 = _io_lu_out_T[15:0]; // @[AccessMemory.scala 14:41]
  wire [63:0] _io_lu_out_T_7 = {io_lu_out_hi_1,io_lu_out_lo_1}; // @[Cat.scala 30:58]
  wire [31:0] io_lu_out_hi_2 = _io_lu_out_T[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] io_lu_out_lo_2 = _io_lu_out_T[31:0]; // @[AccessMemory.scala 15:41]
  wire [63:0] _io_lu_out_T_11 = {io_lu_out_hi_2,io_lu_out_lo_2}; // @[Cat.scala 30:58]
  wire [63:0] _io_lu_out_T_14 = {56'h0,io_lu_out_lo}; // @[Cat.scala 30:58]
  wire [63:0] _io_lu_out_T_16 = {48'h0,io_lu_out_lo_1}; // @[Cat.scala 30:58]
  wire [63:0] _io_lu_out_T_18 = {32'h0,io_lu_out_lo_2}; // @[Cat.scala 30:58]
  wire [63:0] _io_lu_out_T_20 = 7'h1 == io_lu_code ? _io_lu_out_T_3 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _io_lu_out_T_22 = 7'h2 == io_lu_code ? _io_lu_out_T_7 : _io_lu_out_T_20; // @[Mux.scala 80:57]
  wire [63:0] _io_lu_out_T_24 = 7'h4 == io_lu_code ? _io_lu_out_T_11 : _io_lu_out_T_22; // @[Mux.scala 80:57]
  wire [63:0] _io_lu_out_T_26 = 7'h8 == io_lu_code ? _io_lu_out_T : _io_lu_out_T_24; // @[Mux.scala 80:57]
  wire [63:0] _io_lu_out_T_28 = 7'h10 == io_lu_code ? _io_lu_out_T_14 : _io_lu_out_T_26; // @[Mux.scala 80:57]
  wire [63:0] _io_lu_out_T_30 = 7'h20 == io_lu_code ? _io_lu_out_T_16 : _io_lu_out_T_28; // @[Mux.scala 80:57]
  assign io_lu_out = 7'h40 == io_lu_code ? _io_lu_out_T_18 : _io_lu_out_T_30; // @[Mux.scala 80:57]
endmodule
module WriteBack(
  input  [6:0]  io_fu_code,
  input  [63:0] io_alu_out,
  input  [63:0] io_bu_out,
  input  [63:0] io_mu_out,
  input  [63:0] io_du_out,
  input  [63:0] io_lu_out,
  input  [63:0] io_csru_out,
  output [63:0] io_out
);
  wire [63:0] _io_out_T_1 = 7'h1 == io_fu_code ? io_alu_out : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _io_out_T_3 = 7'h2 == io_fu_code ? io_bu_out : _io_out_T_1; // @[Mux.scala 80:57]
  wire [63:0] _io_out_T_5 = 7'h4 == io_fu_code ? io_lu_out : _io_out_T_3; // @[Mux.scala 80:57]
  wire [63:0] _io_out_T_7 = 7'h8 == io_fu_code ? 64'h0 : _io_out_T_5; // @[Mux.scala 80:57]
  wire [63:0] _io_out_T_9 = 7'h10 == io_fu_code ? io_mu_out : _io_out_T_7; // @[Mux.scala 80:57]
  wire [63:0] _io_out_T_11 = 7'h20 == io_fu_code ? io_du_out : _io_out_T_9; // @[Mux.scala 80:57]
  assign io_out = 7'h40 == io_fu_code ? io_csru_out : _io_out_T_11; // @[Mux.scala 80:57]
endmodule
module Mul(
  input          clock,
  input          reset,
  input          io_en,
  input  [64:0]  io_x,
  input  [64:0]  io_y,
  output [129:0] io_out,
  output         io_stall
);
`ifdef RANDOMIZE_REG_INIT
  reg [159:0] _RAND_0;
  reg [95:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [159:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [129:0] x; // @[Mul.scala 14:20]
  reg [64:0] y; // @[Mul.scala 15:20]
  reg [6:0] cnt; // @[Mul.scala 16:22]
  reg [129:0] sum; // @[Mul.scala 17:22]
  reg [1:0] state; // @[Mul.scala 20:24]
  wire  _T = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_1 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_2 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_1 = cnt == 7'h40 ? 2'h3 : state; // @[Mul.scala 30:31 Mul.scala 30:38 Mul.scala 20:24]
  wire  _T_4 = 2'h3 == state; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_2 = _T_4 ? 2'h0 : state; // @[Conditional.scala 39:67 Mul.scala 33:19 Mul.scala 20:24]
  wire [64:0] x_hi = io_x[64] ? 65'h1ffffffffffffffff : 65'h0; // @[Bitwise.scala 72:12]
  wire [129:0] _x_T_2 = {x_hi,io_x}; // @[Cat.scala 30:58]
  wire [130:0] _x_T_3 = {x, 1'h0}; // @[Mul.scala 44:16]
  wire [64:0] _y_T = {{1'd0}, y[64:1]}; // @[Mul.scala 45:16]
  wire [6:0] _cnt_T_1 = cnt + 7'h1; // @[Mul.scala 46:20]
  wire [129:0] _sum_T_1 = y[0] ? x : 130'h0; // @[Mul.scala 47:25]
  wire [129:0] _sum_T_3 = sum + _sum_T_1; // @[Mul.scala 47:20]
  wire [130:0] _GEN_6 = state == 2'h2 ? _x_T_3 : {{1'd0}, x}; // @[Mul.scala 43:33 Mul.scala 44:11 Mul.scala 14:20]
  wire [130:0] _GEN_10 = state == 2'h1 ? {{1'd0}, _x_T_2} : _GEN_6; // @[Mul.scala 37:26 Mul.scala 38:11]
  assign io_out = sum; // @[Mul.scala 50:12]
  assign io_stall = ~(state == 2'h3 | state == 2'h0 & ~io_en); // @[Mul.scala 51:17]
  always @(posedge clock) begin
    if (reset) begin // @[Mul.scala 14:20]
      x <= 130'h0; // @[Mul.scala 14:20]
    end else begin
      x <= _GEN_10[129:0];
    end
    if (reset) begin // @[Mul.scala 15:20]
      y <= 65'h0; // @[Mul.scala 15:20]
    end else if (state == 2'h1) begin // @[Mul.scala 37:26]
      y <= io_y; // @[Mul.scala 39:11]
    end else if (state == 2'h2) begin // @[Mul.scala 43:33]
      y <= _y_T; // @[Mul.scala 45:11]
    end
    if (reset) begin // @[Mul.scala 16:22]
      cnt <= 7'h0; // @[Mul.scala 16:22]
    end else if (state == 2'h1) begin // @[Mul.scala 37:26]
      cnt <= 7'h0; // @[Mul.scala 40:13]
    end else if (state == 2'h2) begin // @[Mul.scala 43:33]
      cnt <= _cnt_T_1; // @[Mul.scala 46:13]
    end
    if (reset) begin // @[Mul.scala 17:22]
      sum <= 130'h0; // @[Mul.scala 17:22]
    end else if (state == 2'h1) begin // @[Mul.scala 37:26]
      sum <= 130'h0; // @[Mul.scala 41:13]
    end else if (state == 2'h2) begin // @[Mul.scala 43:33]
      sum <= _sum_T_3; // @[Mul.scala 47:13]
    end
    if (reset) begin // @[Mul.scala 20:24]
      state <= 2'h0; // @[Mul.scala 20:24]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_en) begin // @[Mul.scala 24:24]
        state <= 2'h1; // @[Mul.scala 24:31]
      end
    end else if (_T_1) begin // @[Conditional.scala 39:67]
      state <= 2'h2; // @[Mul.scala 27:19]
    end else if (_T_2) begin // @[Conditional.scala 39:67]
      state <= _GEN_1;
    end else begin
      state <= _GEN_2;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {5{`RANDOM}};
  x = _RAND_0[129:0];
  _RAND_1 = {3{`RANDOM}};
  y = _RAND_1[64:0];
  _RAND_2 = {1{`RANDOM}};
  cnt = _RAND_2[6:0];
  _RAND_3 = {5{`RANDOM}};
  sum = _RAND_3[129:0];
  _RAND_4 = {1{`RANDOM}};
  state = _RAND_4[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MU(
  input         clock,
  input         reset,
  input         io_en,
  input  [1:0]  io_mu_code,
  input  [63:0] io_op1,
  input  [63:0] io_op2,
  output [63:0] io_mu_out,
  output [63:0] io_stall
);
  wire  mul_clock; // @[Mul.scala 69:21]
  wire  mul_reset; // @[Mul.scala 69:21]
  wire  mul_io_en; // @[Mul.scala 69:21]
  wire [64:0] mul_io_x; // @[Mul.scala 69:21]
  wire [64:0] mul_io_y; // @[Mul.scala 69:21]
  wire [129:0] mul_io_out; // @[Mul.scala 69:21]
  wire  mul_io_stall; // @[Mul.scala 69:21]
  wire [129:0] _mu_out_T_1 = mul_io_out + 130'h1; // @[Mul.scala 76:36]
  wire [31:0] mu_out_hi = _mu_out_T_1[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] mu_out_lo = _mu_out_T_1[31:0]; // @[Mul.scala 67:41]
  wire [63:0] _mu_out_T_4 = {mu_out_hi,mu_out_lo}; // @[Cat.scala 30:58]
  wire [129:0] _mu_out_T_6 = 2'h1 == io_mu_code ? mul_io_out : 130'h0; // @[Mux.scala 80:57]
  wire [129:0] mu_out = 2'h2 == io_mu_code ? {{66'd0}, _mu_out_T_4} : _mu_out_T_6; // @[Mux.scala 80:57]
  Mul mul ( // @[Mul.scala 69:21]
    .clock(mul_clock),
    .reset(mul_reset),
    .io_en(mul_io_en),
    .io_x(mul_io_x),
    .io_y(mul_io_y),
    .io_out(mul_io_out),
    .io_stall(mul_io_stall)
  );
  assign io_mu_out = mu_out[63:0]; // @[Mul.scala 79:17]
  assign io_stall = {{63'd0}, mul_io_stall}; // @[Mul.scala 80:17]
  assign mul_clock = clock;
  assign mul_reset = reset;
  assign mul_io_en = io_en; // @[Mul.scala 70:17]
  assign mul_io_x = {{1'd0}, io_op1}; // @[Mul.scala 71:17]
  assign mul_io_y = {{1'd0}, io_op2}; // @[Mul.scala 72:17]
endmodule
module CorrelationConflict(
  input        io_rs_valid,
  input        io_rd_valid,
  input        io_rs1_en,
  input        io_rs2_en,
  input  [4:0] io_rs1_addr,
  input  [4:0] io_rs2_addr,
  input        io_rd_en,
  input  [4:0] io_rd_addr,
  output       io_conflict
);
  wire  inst_valid = io_rs_valid & io_rd_valid; // @[PipelineReg.scala 166:39]
  wire  rs1_conflict = io_rs1_en & io_rs1_addr == io_rd_addr; // @[PipelineReg.scala 167:37]
  wire  rs2_conflict = io_rs2_en & io_rs2_addr == io_rd_addr; // @[PipelineReg.scala 168:37]
  wire  rd_valid = io_rd_addr != 5'h0 & io_rd_en; // @[PipelineReg.scala 169:48]
  assign io_conflict = inst_valid & rd_valid & (rs1_conflict | rs2_conflict); // @[PipelineReg.scala 171:43]
endmodule
module RegfileConflict(
  input        io_rs_valid,
  input        io_rs1_en,
  input        io_rs2_en,
  input  [4:0] io_rs1_addr,
  input  [4:0] io_rs2_addr,
  input        io_rd1_valid,
  input        io_rd1_en,
  input  [4:0] io_rd1_addr,
  input        io_rd2_valid,
  input        io_rd2_en,
  input  [4:0] io_rd2_addr,
  input        io_rd3_valid,
  input        io_rd3_en,
  input  [4:0] io_rd3_addr,
  output       io_conflict
);
  wire  cconflict1_io_rs_valid; // @[PipelineReg.scala 194:28]
  wire  cconflict1_io_rd_valid; // @[PipelineReg.scala 194:28]
  wire  cconflict1_io_rs1_en; // @[PipelineReg.scala 194:28]
  wire  cconflict1_io_rs2_en; // @[PipelineReg.scala 194:28]
  wire [4:0] cconflict1_io_rs1_addr; // @[PipelineReg.scala 194:28]
  wire [4:0] cconflict1_io_rs2_addr; // @[PipelineReg.scala 194:28]
  wire  cconflict1_io_rd_en; // @[PipelineReg.scala 194:28]
  wire [4:0] cconflict1_io_rd_addr; // @[PipelineReg.scala 194:28]
  wire  cconflict1_io_conflict; // @[PipelineReg.scala 194:28]
  wire  cconflict2_io_rs_valid; // @[PipelineReg.scala 195:28]
  wire  cconflict2_io_rd_valid; // @[PipelineReg.scala 195:28]
  wire  cconflict2_io_rs1_en; // @[PipelineReg.scala 195:28]
  wire  cconflict2_io_rs2_en; // @[PipelineReg.scala 195:28]
  wire [4:0] cconflict2_io_rs1_addr; // @[PipelineReg.scala 195:28]
  wire [4:0] cconflict2_io_rs2_addr; // @[PipelineReg.scala 195:28]
  wire  cconflict2_io_rd_en; // @[PipelineReg.scala 195:28]
  wire [4:0] cconflict2_io_rd_addr; // @[PipelineReg.scala 195:28]
  wire  cconflict2_io_conflict; // @[PipelineReg.scala 195:28]
  wire  cconflict3_io_rs_valid; // @[PipelineReg.scala 196:28]
  wire  cconflict3_io_rd_valid; // @[PipelineReg.scala 196:28]
  wire  cconflict3_io_rs1_en; // @[PipelineReg.scala 196:28]
  wire  cconflict3_io_rs2_en; // @[PipelineReg.scala 196:28]
  wire [4:0] cconflict3_io_rs1_addr; // @[PipelineReg.scala 196:28]
  wire [4:0] cconflict3_io_rs2_addr; // @[PipelineReg.scala 196:28]
  wire  cconflict3_io_rd_en; // @[PipelineReg.scala 196:28]
  wire [4:0] cconflict3_io_rd_addr; // @[PipelineReg.scala 196:28]
  wire  cconflict3_io_conflict; // @[PipelineReg.scala 196:28]
  CorrelationConflict cconflict1 ( // @[PipelineReg.scala 194:28]
    .io_rs_valid(cconflict1_io_rs_valid),
    .io_rd_valid(cconflict1_io_rd_valid),
    .io_rs1_en(cconflict1_io_rs1_en),
    .io_rs2_en(cconflict1_io_rs2_en),
    .io_rs1_addr(cconflict1_io_rs1_addr),
    .io_rs2_addr(cconflict1_io_rs2_addr),
    .io_rd_en(cconflict1_io_rd_en),
    .io_rd_addr(cconflict1_io_rd_addr),
    .io_conflict(cconflict1_io_conflict)
  );
  CorrelationConflict cconflict2 ( // @[PipelineReg.scala 195:28]
    .io_rs_valid(cconflict2_io_rs_valid),
    .io_rd_valid(cconflict2_io_rd_valid),
    .io_rs1_en(cconflict2_io_rs1_en),
    .io_rs2_en(cconflict2_io_rs2_en),
    .io_rs1_addr(cconflict2_io_rs1_addr),
    .io_rs2_addr(cconflict2_io_rs2_addr),
    .io_rd_en(cconflict2_io_rd_en),
    .io_rd_addr(cconflict2_io_rd_addr),
    .io_conflict(cconflict2_io_conflict)
  );
  CorrelationConflict cconflict3 ( // @[PipelineReg.scala 196:28]
    .io_rs_valid(cconflict3_io_rs_valid),
    .io_rd_valid(cconflict3_io_rd_valid),
    .io_rs1_en(cconflict3_io_rs1_en),
    .io_rs2_en(cconflict3_io_rs2_en),
    .io_rs1_addr(cconflict3_io_rs1_addr),
    .io_rs2_addr(cconflict3_io_rs2_addr),
    .io_rd_en(cconflict3_io_rd_en),
    .io_rd_addr(cconflict3_io_rd_addr),
    .io_conflict(cconflict3_io_conflict)
  );
  assign io_conflict = cconflict1_io_conflict | cconflict2_io_conflict | cconflict3_io_conflict; // @[PipelineReg.scala 225:69]
  assign cconflict1_io_rs_valid = io_rs_valid; // @[PipelineReg.scala 198:29]
  assign cconflict1_io_rd_valid = io_rd1_valid; // @[PipelineReg.scala 199:29]
  assign cconflict1_io_rs1_en = io_rs1_en; // @[PipelineReg.scala 200:29]
  assign cconflict1_io_rs2_en = io_rs2_en; // @[PipelineReg.scala 201:29]
  assign cconflict1_io_rs1_addr = io_rs1_addr; // @[PipelineReg.scala 202:29]
  assign cconflict1_io_rs2_addr = io_rs2_addr; // @[PipelineReg.scala 203:29]
  assign cconflict1_io_rd_en = io_rd1_en; // @[PipelineReg.scala 204:29]
  assign cconflict1_io_rd_addr = io_rd1_addr; // @[PipelineReg.scala 205:29]
  assign cconflict2_io_rs_valid = io_rs_valid; // @[PipelineReg.scala 207:29]
  assign cconflict2_io_rd_valid = io_rd2_valid; // @[PipelineReg.scala 208:29]
  assign cconflict2_io_rs1_en = io_rs1_en; // @[PipelineReg.scala 209:29]
  assign cconflict2_io_rs2_en = io_rs2_en; // @[PipelineReg.scala 210:29]
  assign cconflict2_io_rs1_addr = io_rs1_addr; // @[PipelineReg.scala 211:29]
  assign cconflict2_io_rs2_addr = io_rs2_addr; // @[PipelineReg.scala 212:29]
  assign cconflict2_io_rd_en = io_rd2_en; // @[PipelineReg.scala 213:29]
  assign cconflict2_io_rd_addr = io_rd2_addr; // @[PipelineReg.scala 214:29]
  assign cconflict3_io_rs_valid = io_rs_valid; // @[PipelineReg.scala 216:29]
  assign cconflict3_io_rd_valid = io_rd3_valid; // @[PipelineReg.scala 217:29]
  assign cconflict3_io_rs1_en = io_rs1_en; // @[PipelineReg.scala 218:29]
  assign cconflict3_io_rs2_en = io_rs2_en; // @[PipelineReg.scala 219:29]
  assign cconflict3_io_rs1_addr = io_rs1_addr; // @[PipelineReg.scala 220:29]
  assign cconflict3_io_rs2_addr = io_rs2_addr; // @[PipelineReg.scala 221:29]
  assign cconflict3_io_rd_en = io_rd3_en; // @[PipelineReg.scala 222:29]
  assign cconflict3_io_rd_addr = io_rd3_addr; // @[PipelineReg.scala 223:29]
endmodule
module Fence(
  input   clock,
  input   reset,
  input   io_go,
  output  io_ok,
  output  io_ifence_req,
  input   io_ifence_done,
  output  io_dfence_req,
  input   io_dfence_done
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[Fence.scala 19:24]
  wire  _T = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_1 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_2 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_1 = io_dfence_done ? 3'h3 : state; // @[Fence.scala 29:33 Fence.scala 29:40 Fence.scala 19:24]
  wire  _T_3 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_2 = io_ifence_done ? 3'h4 : state; // @[Fence.scala 32:33 Fence.scala 32:40 Fence.scala 19:24]
  wire  _T_4 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_3 = _T_4 ? 3'h0 : state; // @[Conditional.scala 39:67 Fence.scala 35:19 Fence.scala 19:24]
  wire [2:0] _GEN_4 = _T_3 ? _GEN_2 : _GEN_3; // @[Conditional.scala 39:67]
  assign io_ok = state == 3'h0 & ~io_go | state == 3'h4 | state == 3'h1; // @[Fence.scala 39:70]
  assign io_ifence_req = state == 3'h3; // @[Fence.scala 41:28]
  assign io_dfence_req = state == 3'h2; // @[Fence.scala 40:28]
  always @(posedge clock) begin
    if (reset) begin // @[Fence.scala 19:24]
      state <= 3'h0; // @[Fence.scala 19:24]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_go) begin // @[Fence.scala 23:24]
        state <= 3'h1; // @[Fence.scala 23:31]
      end
    end else if (_T_1) begin // @[Conditional.scala 39:67]
      state <= 3'h2; // @[Fence.scala 26:19]
    end else if (_T_2) begin // @[Conditional.scala 39:67]
      state <= _GEN_1;
    end else begin
      state <= _GEN_4;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IDReg(
  input         clock,
  input         reset,
  input         io_en,
  input         io_in_valid,
  input  [63:0] io_in_pc,
  output        io_out_valid,
  output [63:0] io_out_pc,
  output [63:0] io_imem__addr,
  output        io_imem__en,
  input  [31:0] io_imem__data,
  output [31:0] io_inst
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  valid; // @[Reg.scala 27:20]
  reg [63:0] pc; // @[Reg.scala 27:20]
  assign io_out_valid = valid; // @[PipelineReg.scala 31:21]
  assign io_out_pc = pc; // @[PipelineReg.scala 32:21]
  assign io_imem__addr = io_in_pc; // @[PipelineReg.scala 26:21]
  assign io_imem__en = io_en; // @[PipelineReg.scala 27:21]
  assign io_inst = io_imem__data; // @[PipelineReg.scala 28:21]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 27:20]
      valid <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      valid <= io_in_valid; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      pc <= 64'h7ffffffc; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      pc <= io_in_pc; // @[Reg.scala 28:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  pc = _RAND_1[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ExeReg(
  input         clock,
  input         reset,
  input         io_en,
  input         io_in_valid,
  input  [63:0] io_in_pc,
  input  [31:0] io_in_inst,
  input         io_in_rd_en,
  input  [4:0]  io_in_rd_addr,
  input  [63:0] io_in_imm,
  input  [63:0] io_in_op1,
  input  [63:0] io_in_op2,
  input  [6:0]  io_in_fu_code,
  input  [15:0] io_in_alu_code,
  input  [7:0]  io_in_bu_code,
  input  [6:0]  io_in_lu_code,
  input  [3:0]  io_in_su_code,
  input  [1:0]  io_in_mu_code,
  input  [7:0]  io_in_du_code,
  input  [7:0]  io_in_csru_code,
  input  [4:0]  io_in_rs1_addr,
  input         io_in_putch,
  output        io_out_valid,
  output [63:0] io_out_pc,
  output [31:0] io_out_inst,
  output        io_out_rd_en,
  output [4:0]  io_out_rd_addr,
  output [63:0] io_out_imm,
  output [63:0] io_out_op1,
  output [63:0] io_out_op2,
  output [6:0]  io_out_fu_code,
  output [15:0] io_out_alu_code,
  output [7:0]  io_out_bu_code,
  output [6:0]  io_out_lu_code,
  output [3:0]  io_out_su_code,
  output [1:0]  io_out_mu_code,
  output [7:0]  io_out_du_code,
  output [7:0]  io_out_csru_code,
  output [4:0]  io_out_rs1_addr,
  output        io_out_putch
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  reg  reg_valid; // @[Reg.scala 27:20]
  reg [63:0] reg_pc; // @[Reg.scala 27:20]
  reg [31:0] reg_inst; // @[Reg.scala 27:20]
  reg  reg_rd_en; // @[Reg.scala 27:20]
  reg [4:0] reg_rd_addr; // @[Reg.scala 27:20]
  reg [63:0] reg_imm; // @[Reg.scala 27:20]
  reg [63:0] reg_op1; // @[Reg.scala 27:20]
  reg [63:0] reg_op2; // @[Reg.scala 27:20]
  reg [6:0] reg_fu_code; // @[Reg.scala 27:20]
  reg [15:0] reg_alu_code; // @[Reg.scala 27:20]
  reg [7:0] reg_bu_code; // @[Reg.scala 27:20]
  reg [6:0] reg_lu_code; // @[Reg.scala 27:20]
  reg [3:0] reg_su_code; // @[Reg.scala 27:20]
  reg [1:0] reg_mu_code; // @[Reg.scala 27:20]
  reg [7:0] reg_du_code; // @[Reg.scala 27:20]
  reg [7:0] reg_csru_code; // @[Reg.scala 27:20]
  reg [4:0] reg_rs1_addr; // @[Reg.scala 27:20]
  reg  reg_putch; // @[Reg.scala 27:20]
  assign io_out_valid = reg_valid; // @[PipelineReg.scala 66:10]
  assign io_out_pc = reg_pc; // @[PipelineReg.scala 66:10]
  assign io_out_inst = reg_inst; // @[PipelineReg.scala 66:10]
  assign io_out_rd_en = reg_rd_en; // @[PipelineReg.scala 66:10]
  assign io_out_rd_addr = reg_rd_addr; // @[PipelineReg.scala 66:10]
  assign io_out_imm = reg_imm; // @[PipelineReg.scala 66:10]
  assign io_out_op1 = reg_op1; // @[PipelineReg.scala 66:10]
  assign io_out_op2 = reg_op2; // @[PipelineReg.scala 66:10]
  assign io_out_fu_code = reg_fu_code; // @[PipelineReg.scala 66:10]
  assign io_out_alu_code = reg_alu_code; // @[PipelineReg.scala 66:10]
  assign io_out_bu_code = reg_bu_code; // @[PipelineReg.scala 66:10]
  assign io_out_lu_code = reg_lu_code; // @[PipelineReg.scala 66:10]
  assign io_out_su_code = reg_su_code; // @[PipelineReg.scala 66:10]
  assign io_out_mu_code = reg_mu_code; // @[PipelineReg.scala 66:10]
  assign io_out_du_code = reg_du_code; // @[PipelineReg.scala 66:10]
  assign io_out_csru_code = reg_csru_code; // @[PipelineReg.scala 66:10]
  assign io_out_rs1_addr = reg_rs1_addr; // @[PipelineReg.scala 66:10]
  assign io_out_putch = reg_putch; // @[PipelineReg.scala 66:10]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 27:20]
      reg_valid <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_valid <= io_in_valid; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_pc <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_pc <= io_in_pc; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_inst <= 32'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_inst <= io_in_inst; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_rd_en <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_rd_en <= io_in_rd_en; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_rd_addr <= 5'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_rd_addr <= io_in_rd_addr; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_imm <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_imm <= io_in_imm; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_op1 <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_op1 <= io_in_op1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_op2 <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_op2 <= io_in_op2; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_fu_code <= 7'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_fu_code <= io_in_fu_code; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_alu_code <= 16'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_alu_code <= io_in_alu_code; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_bu_code <= 8'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_bu_code <= io_in_bu_code; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_lu_code <= 7'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_lu_code <= io_in_lu_code; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_su_code <= 4'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_su_code <= io_in_su_code; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_mu_code <= 2'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_mu_code <= io_in_mu_code; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_du_code <= 8'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_du_code <= io_in_du_code; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_csru_code <= 8'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_csru_code <= io_in_csru_code; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_rs1_addr <= 5'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_rs1_addr <= io_in_rs1_addr; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_putch <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_putch <= io_in_putch; // @[Reg.scala 28:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_valid = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  reg_pc = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  reg_inst = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  reg_rd_en = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  reg_rd_addr = _RAND_4[4:0];
  _RAND_5 = {2{`RANDOM}};
  reg_imm = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  reg_op1 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  reg_op2 = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  reg_fu_code = _RAND_8[6:0];
  _RAND_9 = {1{`RANDOM}};
  reg_alu_code = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  reg_bu_code = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  reg_lu_code = _RAND_11[6:0];
  _RAND_12 = {1{`RANDOM}};
  reg_su_code = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  reg_mu_code = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  reg_du_code = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  reg_csru_code = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  reg_rs1_addr = _RAND_16[4:0];
  _RAND_17 = {1{`RANDOM}};
  reg_putch = _RAND_17[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MemReg(
  input         clock,
  input         reset,
  input         io_en,
  input         io_in_valid,
  input  [63:0] io_in_pc,
  input  [31:0] io_in_inst,
  input         io_in_rd_en,
  input  [4:0]  io_in_rd_addr,
  input  [63:0] io_in_imm,
  input  [63:0] io_in_op1,
  input  [63:0] io_in_op2,
  input  [63:0] io_in_alu_out,
  input  [63:0] io_in_bu_out,
  input  [63:0] io_in_mu_out,
  input  [63:0] io_in_du_out,
  input  [63:0] io_in_csru_out,
  input  [6:0]  io_in_fu_code,
  input  [6:0]  io_in_lu_code,
  input  [3:0]  io_in_su_code,
  input         io_in_putch,
  input         io_in_csr_wen,
  input  [11:0] io_in_csr_waddr,
  input  [63:0] io_in_csr_wdata,
  output        io_out_valid,
  output [63:0] io_out_pc,
  output [31:0] io_out_inst,
  output        io_out_rd_en,
  output [4:0]  io_out_rd_addr,
  output [63:0] io_out_imm,
  output [63:0] io_out_op1,
  output [63:0] io_out_op2,
  output [63:0] io_out_alu_out,
  output [63:0] io_out_bu_out,
  output [63:0] io_out_mu_out,
  output [63:0] io_out_du_out,
  output [63:0] io_out_csru_out,
  output [6:0]  io_out_fu_code,
  output [6:0]  io_out_lu_code,
  output [3:0]  io_out_su_code,
  output        io_out_putch,
  output        io_out_csr_wen,
  output [11:0] io_out_csr_waddr,
  output [63:0] io_out_csr_wdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [63:0] _RAND_19;
`endif // RANDOMIZE_REG_INIT
  reg  reg_valid; // @[Reg.scala 27:20]
  reg [63:0] reg_pc; // @[Reg.scala 27:20]
  reg [31:0] reg_inst; // @[Reg.scala 27:20]
  reg  reg_rd_en; // @[Reg.scala 27:20]
  reg [4:0] reg_rd_addr; // @[Reg.scala 27:20]
  reg [63:0] reg_imm; // @[Reg.scala 27:20]
  reg [63:0] reg_op1; // @[Reg.scala 27:20]
  reg [63:0] reg_op2; // @[Reg.scala 27:20]
  reg [63:0] reg_alu_out; // @[Reg.scala 27:20]
  reg [63:0] reg_bu_out; // @[Reg.scala 27:20]
  reg [63:0] reg_mu_out; // @[Reg.scala 27:20]
  reg [63:0] reg_du_out; // @[Reg.scala 27:20]
  reg [63:0] reg_csru_out; // @[Reg.scala 27:20]
  reg [6:0] reg_fu_code; // @[Reg.scala 27:20]
  reg [6:0] reg_lu_code; // @[Reg.scala 27:20]
  reg [3:0] reg_su_code; // @[Reg.scala 27:20]
  reg  reg_putch; // @[Reg.scala 27:20]
  reg  reg_csr_wen; // @[Reg.scala 27:20]
  reg [11:0] reg_csr_waddr; // @[Reg.scala 27:20]
  reg [63:0] reg_csr_wdata; // @[Reg.scala 27:20]
  assign io_out_valid = reg_valid; // @[PipelineReg.scala 110:10]
  assign io_out_pc = reg_pc; // @[PipelineReg.scala 110:10]
  assign io_out_inst = reg_inst; // @[PipelineReg.scala 110:10]
  assign io_out_rd_en = reg_rd_en; // @[PipelineReg.scala 110:10]
  assign io_out_rd_addr = reg_rd_addr; // @[PipelineReg.scala 110:10]
  assign io_out_imm = reg_imm; // @[PipelineReg.scala 110:10]
  assign io_out_op1 = reg_op1; // @[PipelineReg.scala 110:10]
  assign io_out_op2 = reg_op2; // @[PipelineReg.scala 110:10]
  assign io_out_alu_out = reg_alu_out; // @[PipelineReg.scala 110:10]
  assign io_out_bu_out = reg_bu_out; // @[PipelineReg.scala 110:10]
  assign io_out_mu_out = reg_mu_out; // @[PipelineReg.scala 110:10]
  assign io_out_du_out = reg_du_out; // @[PipelineReg.scala 110:10]
  assign io_out_csru_out = reg_csru_out; // @[PipelineReg.scala 110:10]
  assign io_out_fu_code = reg_fu_code; // @[PipelineReg.scala 110:10]
  assign io_out_lu_code = reg_lu_code; // @[PipelineReg.scala 110:10]
  assign io_out_su_code = reg_su_code; // @[PipelineReg.scala 110:10]
  assign io_out_putch = reg_putch; // @[PipelineReg.scala 110:10]
  assign io_out_csr_wen = reg_csr_wen; // @[PipelineReg.scala 110:10]
  assign io_out_csr_waddr = reg_csr_waddr; // @[PipelineReg.scala 110:10]
  assign io_out_csr_wdata = reg_csr_wdata; // @[PipelineReg.scala 110:10]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 27:20]
      reg_valid <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_valid <= io_in_valid; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_pc <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_pc <= io_in_pc; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_inst <= 32'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_inst <= io_in_inst; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_rd_en <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_rd_en <= io_in_rd_en; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_rd_addr <= 5'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_rd_addr <= io_in_rd_addr; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_imm <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_imm <= io_in_imm; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_op1 <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_op1 <= io_in_op1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_op2 <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_op2 <= io_in_op2; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_alu_out <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_alu_out <= io_in_alu_out; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_bu_out <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_bu_out <= io_in_bu_out; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_mu_out <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_mu_out <= io_in_mu_out; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_du_out <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_du_out <= io_in_du_out; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_csru_out <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_csru_out <= io_in_csru_out; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_fu_code <= 7'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_fu_code <= io_in_fu_code; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_lu_code <= 7'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_lu_code <= io_in_lu_code; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_su_code <= 4'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_su_code <= io_in_su_code; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_putch <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_putch <= io_in_putch; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_csr_wen <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_csr_wen <= io_in_csr_wen; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_csr_waddr <= 12'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_csr_waddr <= io_in_csr_waddr; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_csr_wdata <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_csr_wdata <= io_in_csr_wdata; // @[Reg.scala 28:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_valid = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  reg_pc = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  reg_inst = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  reg_rd_en = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  reg_rd_addr = _RAND_4[4:0];
  _RAND_5 = {2{`RANDOM}};
  reg_imm = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  reg_op1 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  reg_op2 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  reg_alu_out = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  reg_bu_out = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  reg_mu_out = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  reg_du_out = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  reg_csru_out = _RAND_12[63:0];
  _RAND_13 = {1{`RANDOM}};
  reg_fu_code = _RAND_13[6:0];
  _RAND_14 = {1{`RANDOM}};
  reg_lu_code = _RAND_14[6:0];
  _RAND_15 = {1{`RANDOM}};
  reg_su_code = _RAND_15[3:0];
  _RAND_16 = {1{`RANDOM}};
  reg_putch = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  reg_csr_wen = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  reg_csr_waddr = _RAND_18[11:0];
  _RAND_19 = {2{`RANDOM}};
  reg_csr_wdata = _RAND_19[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module WBReg(
  input         clock,
  input         reset,
  input         io_en,
  input         io_in_valid,
  input  [63:0] io_in_pc,
  input  [31:0] io_in_inst,
  input         io_in_rd_en,
  input  [4:0]  io_in_rd_addr,
  input  [63:0] io_in_alu_out,
  input  [63:0] io_in_bu_out,
  input  [63:0] io_in_mu_out,
  input  [63:0] io_in_du_out,
  input  [63:0] io_in_csru_out,
  input  [6:0]  io_in_fu_code,
  input  [6:0]  io_in_lu_code,
  input  [5:0]  io_in_lu_shift,
  input         io_in_putch,
  input         io_in_csr_wen,
  input  [11:0] io_in_csr_waddr,
  input  [63:0] io_in_csr_wdata,
  input         io_in_csr_set_mtip,
  input         io_in_csr_clear_mtip,
  output        io_out_valid,
  output [63:0] io_out_pc,
  output [31:0] io_out_inst,
  output        io_out_rd_en,
  output [4:0]  io_out_rd_addr,
  output [63:0] io_out_alu_out,
  output [63:0] io_out_bu_out,
  output [63:0] io_out_mu_out,
  output [63:0] io_out_du_out,
  output [63:0] io_out_csru_out,
  output [6:0]  io_out_fu_code,
  output [6:0]  io_out_lu_code,
  output [5:0]  io_out_lu_shift,
  output        io_out_putch,
  output        io_out_csr_wen,
  output [11:0] io_out_csr_waddr,
  output [63:0] io_out_csr_wdata,
  output        io_out_csr_set_mtip,
  output        io_out_csr_clear_mtip
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  reg  reg_valid; // @[Reg.scala 27:20]
  reg [63:0] reg_pc; // @[Reg.scala 27:20]
  reg [31:0] reg_inst; // @[Reg.scala 27:20]
  reg  reg_rd_en; // @[Reg.scala 27:20]
  reg [4:0] reg_rd_addr; // @[Reg.scala 27:20]
  reg [63:0] reg_alu_out; // @[Reg.scala 27:20]
  reg [63:0] reg_bu_out; // @[Reg.scala 27:20]
  reg [63:0] reg_mu_out; // @[Reg.scala 27:20]
  reg [63:0] reg_du_out; // @[Reg.scala 27:20]
  reg [63:0] reg_csru_out; // @[Reg.scala 27:20]
  reg [6:0] reg_fu_code; // @[Reg.scala 27:20]
  reg [6:0] reg_lu_code; // @[Reg.scala 27:20]
  reg [5:0] reg_lu_shift; // @[Reg.scala 27:20]
  reg  reg_putch; // @[Reg.scala 27:20]
  reg  reg_csr_wen; // @[Reg.scala 27:20]
  reg [11:0] reg_csr_waddr; // @[Reg.scala 27:20]
  reg [63:0] reg_csr_wdata; // @[Reg.scala 27:20]
  reg  reg_csr_set_mtip; // @[Reg.scala 27:20]
  reg  reg_csr_clear_mtip; // @[Reg.scala 27:20]
  assign io_out_valid = reg_valid; // @[PipelineReg.scala 150:10]
  assign io_out_pc = reg_pc; // @[PipelineReg.scala 150:10]
  assign io_out_inst = reg_inst; // @[PipelineReg.scala 150:10]
  assign io_out_rd_en = reg_rd_en; // @[PipelineReg.scala 150:10]
  assign io_out_rd_addr = reg_rd_addr; // @[PipelineReg.scala 150:10]
  assign io_out_alu_out = reg_alu_out; // @[PipelineReg.scala 150:10]
  assign io_out_bu_out = reg_bu_out; // @[PipelineReg.scala 150:10]
  assign io_out_mu_out = reg_mu_out; // @[PipelineReg.scala 150:10]
  assign io_out_du_out = reg_du_out; // @[PipelineReg.scala 150:10]
  assign io_out_csru_out = reg_csru_out; // @[PipelineReg.scala 150:10]
  assign io_out_fu_code = reg_fu_code; // @[PipelineReg.scala 150:10]
  assign io_out_lu_code = reg_lu_code; // @[PipelineReg.scala 150:10]
  assign io_out_lu_shift = reg_lu_shift; // @[PipelineReg.scala 150:10]
  assign io_out_putch = reg_putch; // @[PipelineReg.scala 150:10]
  assign io_out_csr_wen = reg_csr_wen; // @[PipelineReg.scala 150:10]
  assign io_out_csr_waddr = reg_csr_waddr; // @[PipelineReg.scala 150:10]
  assign io_out_csr_wdata = reg_csr_wdata; // @[PipelineReg.scala 150:10]
  assign io_out_csr_set_mtip = reg_csr_set_mtip; // @[PipelineReg.scala 150:10]
  assign io_out_csr_clear_mtip = reg_csr_clear_mtip; // @[PipelineReg.scala 150:10]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 27:20]
      reg_valid <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_valid <= io_in_valid; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_pc <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_pc <= io_in_pc; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_inst <= 32'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_inst <= io_in_inst; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_rd_en <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_rd_en <= io_in_rd_en; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_rd_addr <= 5'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_rd_addr <= io_in_rd_addr; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_alu_out <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_alu_out <= io_in_alu_out; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_bu_out <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_bu_out <= io_in_bu_out; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_mu_out <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_mu_out <= io_in_mu_out; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_du_out <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_du_out <= io_in_du_out; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_csru_out <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_csru_out <= io_in_csru_out; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_fu_code <= 7'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_fu_code <= io_in_fu_code; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_lu_code <= 7'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_lu_code <= io_in_lu_code; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_lu_shift <= 6'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_lu_shift <= io_in_lu_shift; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_putch <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_putch <= io_in_putch; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_csr_wen <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_csr_wen <= io_in_csr_wen; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_csr_waddr <= 12'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_csr_waddr <= io_in_csr_waddr; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_csr_wdata <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_csr_wdata <= io_in_csr_wdata; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_csr_set_mtip <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_csr_set_mtip <= io_in_csr_set_mtip; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_csr_clear_mtip <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_en) begin // @[Reg.scala 28:19]
      reg_csr_clear_mtip <= io_in_csr_clear_mtip; // @[Reg.scala 28:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_valid = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  reg_pc = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  reg_inst = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  reg_rd_en = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  reg_rd_addr = _RAND_4[4:0];
  _RAND_5 = {2{`RANDOM}};
  reg_alu_out = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  reg_bu_out = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  reg_mu_out = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  reg_du_out = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  reg_csru_out = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  reg_fu_code = _RAND_10[6:0];
  _RAND_11 = {1{`RANDOM}};
  reg_lu_code = _RAND_11[6:0];
  _RAND_12 = {1{`RANDOM}};
  reg_lu_shift = _RAND_12[5:0];
  _RAND_13 = {1{`RANDOM}};
  reg_putch = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  reg_csr_wen = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  reg_csr_waddr = _RAND_15[11:0];
  _RAND_16 = {2{`RANDOM}};
  reg_csr_wdata = _RAND_16[63:0];
  _RAND_17 = {1{`RANDOM}};
  reg_csr_set_mtip = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  reg_csr_clear_mtip = _RAND_18[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Core(
  input         clock,
  input         reset,
  output [63:0] io_imem_addr,
  output        io_imem_en,
  input  [31:0] io_imem_data,
  input         io_imem_ok,
  output        io_dmem_en,
  output        io_dmem_op,
  output [63:0] io_dmem_addr,
  output [63:0] io_dmem_wdata,
  output [7:0]  io_dmem_wmask,
  output [31:0] io_dmem_transfer,
  input         io_dmem_ok,
  input  [63:0] io_dmem_rdata,
  input         io_set_mtip,
  input         io_clear_mtip,
  output        io_ifence_req,
  input         io_ifence_done,
  output        io_dfence_req,
  input         io_dfence_done
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
`endif // RANDOMIZE_REG_INIT
  wire  ifu_reset; // @[Core.scala 19:23]
  wire  ifu_io_jump_en; // @[Core.scala 19:23]
  wire [63:0] ifu_io_jump_pc; // @[Core.scala 19:23]
  wire [63:0] ifu_io_pc; // @[Core.scala 19:23]
  wire [63:0] ifu_io_next_pc; // @[Core.scala 19:23]
  wire  ifu_io_valid; // @[Core.scala 19:23]
  wire [63:0] idu_io_pc; // @[Core.scala 20:23]
  wire [31:0] idu_io_inst; // @[Core.scala 20:23]
  wire  idu_io_rs1_en; // @[Core.scala 20:23]
  wire  idu_io_rs2_en; // @[Core.scala 20:23]
  wire [4:0] idu_io_rs1_addr; // @[Core.scala 20:23]
  wire [4:0] idu_io_rs2_addr; // @[Core.scala 20:23]
  wire [63:0] idu_io_rs1_data; // @[Core.scala 20:23]
  wire [63:0] idu_io_rs2_data; // @[Core.scala 20:23]
  wire  idu_io_rd_en; // @[Core.scala 20:23]
  wire [4:0] idu_io_rd_addr; // @[Core.scala 20:23]
  wire [6:0] idu_io_decode_info_fu_code; // @[Core.scala 20:23]
  wire [15:0] idu_io_decode_info_alu_code; // @[Core.scala 20:23]
  wire [7:0] idu_io_decode_info_bu_code; // @[Core.scala 20:23]
  wire [6:0] idu_io_decode_info_lu_code; // @[Core.scala 20:23]
  wire [3:0] idu_io_decode_info_su_code; // @[Core.scala 20:23]
  wire [1:0] idu_io_decode_info_mu_code; // @[Core.scala 20:23]
  wire [7:0] idu_io_decode_info_du_code; // @[Core.scala 20:23]
  wire [7:0] idu_io_decode_info_csru_code; // @[Core.scala 20:23]
  wire  idu_io_jump_en; // @[Core.scala 20:23]
  wire [63:0] idu_io_jump_pc; // @[Core.scala 20:23]
  wire [63:0] idu_io_op1; // @[Core.scala 20:23]
  wire [63:0] idu_io_op2; // @[Core.scala 20:23]
  wire [63:0] idu_io_imm; // @[Core.scala 20:23]
  wire  idu_io_putch; // @[Core.scala 20:23]
  wire [63:0] idu_io_mtvec; // @[Core.scala 20:23]
  wire [63:0] idu_io_mepc; // @[Core.scala 20:23]
  wire [15:0] ieu_io_alu_code; // @[Core.scala 21:23]
  wire [7:0] ieu_io_bu_code; // @[Core.scala 21:23]
  wire [7:0] ieu_io_du_code; // @[Core.scala 21:23]
  wire [7:0] ieu_io_csru_code; // @[Core.scala 21:23]
  wire [63:0] ieu_io_op1; // @[Core.scala 21:23]
  wire [63:0] ieu_io_op2; // @[Core.scala 21:23]
  wire [63:0] ieu_io_pc; // @[Core.scala 21:23]
  wire [63:0] ieu_io_alu_out; // @[Core.scala 21:23]
  wire [63:0] ieu_io_bu_out; // @[Core.scala 21:23]
  wire [63:0] ieu_io_du_out; // @[Core.scala 21:23]
  wire [63:0] ieu_io_csru_out; // @[Core.scala 21:23]
  wire [4:0] ieu_io_rs1_addr; // @[Core.scala 21:23]
  wire [11:0] ieu_io_csr_raddr; // @[Core.scala 21:23]
  wire [63:0] ieu_io_csr_rdata; // @[Core.scala 21:23]
  wire  ieu_io_csr_wen; // @[Core.scala 21:23]
  wire [11:0] ieu_io_csr_waddr; // @[Core.scala 21:23]
  wire [63:0] ieu_io_csr_wdata; // @[Core.scala 21:23]
  wire  rfu_clock; // @[Core.scala 22:23]
  wire  rfu_reset; // @[Core.scala 22:23]
  wire [4:0] rfu_io_rs1_addr; // @[Core.scala 22:23]
  wire [4:0] rfu_io_rs2_addr; // @[Core.scala 22:23]
  wire [63:0] rfu_io_rs1_data; // @[Core.scala 22:23]
  wire [63:0] rfu_io_rs2_data; // @[Core.scala 22:23]
  wire [4:0] rfu_io_rd_addr; // @[Core.scala 22:23]
  wire [63:0] rfu_io_rd_data; // @[Core.scala 22:23]
  wire  rfu_io_rd_en; // @[Core.scala 22:23]
  wire [63:0] rfu_rf_10; // @[Core.scala 22:23]
  wire  csru_clock; // @[Core.scala 23:23]
  wire  csru_reset; // @[Core.scala 23:23]
  wire [11:0] csru_io_raddr; // @[Core.scala 23:23]
  wire [63:0] csru_io_rdata; // @[Core.scala 23:23]
  wire  csru_io_wen; // @[Core.scala 23:23]
  wire [11:0] csru_io_waddr; // @[Core.scala 23:23]
  wire [63:0] csru_io_wdata; // @[Core.scala 23:23]
  wire  csru_io_set_mtip; // @[Core.scala 23:23]
  wire  csru_io_clear_mtip; // @[Core.scala 23:23]
  wire  csru_io_exception; // @[Core.scala 23:23]
  wire [63:0] csru_io_cause; // @[Core.scala 23:23]
  wire  csru_io_mret; // @[Core.scala 23:23]
  wire [63:0] csru_io_pc; // @[Core.scala 23:23]
  wire [63:0] csru_io_mtvec; // @[Core.scala 23:23]
  wire [63:0] csru_io_mepc; // @[Core.scala 23:23]
  wire  csru_io_time_intr; // @[Core.scala 23:23]
  wire [6:0] preamu_io_lu_code; // @[Core.scala 24:23]
  wire [3:0] preamu_io_su_code; // @[Core.scala 24:23]
  wire [63:0] preamu_io_op1; // @[Core.scala 24:23]
  wire [63:0] preamu_io_op2; // @[Core.scala 24:23]
  wire [63:0] preamu_io_imm; // @[Core.scala 24:23]
  wire [5:0] preamu_io_lu_shift; // @[Core.scala 24:23]
  wire  preamu_io_ren; // @[Core.scala 24:23]
  wire [63:0] preamu_io_raddr; // @[Core.scala 24:23]
  wire  preamu_io_wen; // @[Core.scala 24:23]
  wire [63:0] preamu_io_waddr; // @[Core.scala 24:23]
  wire [63:0] preamu_io_wdata; // @[Core.scala 24:23]
  wire [7:0] preamu_io_wmask; // @[Core.scala 24:23]
  wire [2:0] preamu_io_transfer; // @[Core.scala 24:23]
  wire [6:0] amu_io_lu_code; // @[Core.scala 25:23]
  wire [5:0] amu_io_lu_shift; // @[Core.scala 25:23]
  wire [63:0] amu_io_rdata; // @[Core.scala 25:23]
  wire [63:0] amu_io_lu_out; // @[Core.scala 25:23]
  wire [6:0] wbu_io_fu_code; // @[Core.scala 26:23]
  wire [63:0] wbu_io_alu_out; // @[Core.scala 26:23]
  wire [63:0] wbu_io_bu_out; // @[Core.scala 26:23]
  wire [63:0] wbu_io_mu_out; // @[Core.scala 26:23]
  wire [63:0] wbu_io_du_out; // @[Core.scala 26:23]
  wire [63:0] wbu_io_lu_out; // @[Core.scala 26:23]
  wire [63:0] wbu_io_csru_out; // @[Core.scala 26:23]
  wire [63:0] wbu_io_out; // @[Core.scala 26:23]
  wire  mu_clock; // @[Core.scala 28:23]
  wire  mu_reset; // @[Core.scala 28:23]
  wire  mu_io_en; // @[Core.scala 28:23]
  wire [1:0] mu_io_mu_code; // @[Core.scala 28:23]
  wire [63:0] mu_io_op1; // @[Core.scala 28:23]
  wire [63:0] mu_io_op2; // @[Core.scala 28:23]
  wire [63:0] mu_io_mu_out; // @[Core.scala 28:23]
  wire [63:0] mu_io_stall; // @[Core.scala 28:23]
  wire  rfconflict_io_rs_valid; // @[Core.scala 30:27]
  wire  rfconflict_io_rs1_en; // @[Core.scala 30:27]
  wire  rfconflict_io_rs2_en; // @[Core.scala 30:27]
  wire [4:0] rfconflict_io_rs1_addr; // @[Core.scala 30:27]
  wire [4:0] rfconflict_io_rs2_addr; // @[Core.scala 30:27]
  wire  rfconflict_io_rd1_valid; // @[Core.scala 30:27]
  wire  rfconflict_io_rd1_en; // @[Core.scala 30:27]
  wire [4:0] rfconflict_io_rd1_addr; // @[Core.scala 30:27]
  wire  rfconflict_io_rd2_valid; // @[Core.scala 30:27]
  wire  rfconflict_io_rd2_en; // @[Core.scala 30:27]
  wire [4:0] rfconflict_io_rd2_addr; // @[Core.scala 30:27]
  wire  rfconflict_io_rd3_valid; // @[Core.scala 30:27]
  wire  rfconflict_io_rd3_en; // @[Core.scala 30:27]
  wire [4:0] rfconflict_io_rd3_addr; // @[Core.scala 30:27]
  wire  rfconflict_io_conflict; // @[Core.scala 30:27]
  wire  fence_clock; // @[Core.scala 31:21]
  wire  fence_reset; // @[Core.scala 31:21]
  wire  fence_io_go; // @[Core.scala 31:21]
  wire  fence_io_ok; // @[Core.scala 31:21]
  wire  fence_io_ifence_req; // @[Core.scala 31:21]
  wire  fence_io_ifence_done; // @[Core.scala 31:21]
  wire  fence_io_dfence_req; // @[Core.scala 31:21]
  wire  fence_io_dfence_done; // @[Core.scala 31:21]
  wire  idreg_clock; // @[Core.scala 33:23]
  wire  idreg_reset; // @[Core.scala 33:23]
  wire  idreg_io_en; // @[Core.scala 33:23]
  wire  idreg_io_in_valid; // @[Core.scala 33:23]
  wire [63:0] idreg_io_in_pc; // @[Core.scala 33:23]
  wire  idreg_io_out_valid; // @[Core.scala 33:23]
  wire [63:0] idreg_io_out_pc; // @[Core.scala 33:23]
  wire [63:0] idreg_io_imem__addr; // @[Core.scala 33:23]
  wire  idreg_io_imem__en; // @[Core.scala 33:23]
  wire [31:0] idreg_io_imem__data; // @[Core.scala 33:23]
  wire [31:0] idreg_io_inst; // @[Core.scala 33:23]
  wire  exereg_clock; // @[Core.scala 34:23]
  wire  exereg_reset; // @[Core.scala 34:23]
  wire  exereg_io_en; // @[Core.scala 34:23]
  wire  exereg_io_in_valid; // @[Core.scala 34:23]
  wire [63:0] exereg_io_in_pc; // @[Core.scala 34:23]
  wire [31:0] exereg_io_in_inst; // @[Core.scala 34:23]
  wire  exereg_io_in_rd_en; // @[Core.scala 34:23]
  wire [4:0] exereg_io_in_rd_addr; // @[Core.scala 34:23]
  wire [63:0] exereg_io_in_imm; // @[Core.scala 34:23]
  wire [63:0] exereg_io_in_op1; // @[Core.scala 34:23]
  wire [63:0] exereg_io_in_op2; // @[Core.scala 34:23]
  wire [6:0] exereg_io_in_fu_code; // @[Core.scala 34:23]
  wire [15:0] exereg_io_in_alu_code; // @[Core.scala 34:23]
  wire [7:0] exereg_io_in_bu_code; // @[Core.scala 34:23]
  wire [6:0] exereg_io_in_lu_code; // @[Core.scala 34:23]
  wire [3:0] exereg_io_in_su_code; // @[Core.scala 34:23]
  wire [1:0] exereg_io_in_mu_code; // @[Core.scala 34:23]
  wire [7:0] exereg_io_in_du_code; // @[Core.scala 34:23]
  wire [7:0] exereg_io_in_csru_code; // @[Core.scala 34:23]
  wire [4:0] exereg_io_in_rs1_addr; // @[Core.scala 34:23]
  wire  exereg_io_in_putch; // @[Core.scala 34:23]
  wire  exereg_io_out_valid; // @[Core.scala 34:23]
  wire [63:0] exereg_io_out_pc; // @[Core.scala 34:23]
  wire [31:0] exereg_io_out_inst; // @[Core.scala 34:23]
  wire  exereg_io_out_rd_en; // @[Core.scala 34:23]
  wire [4:0] exereg_io_out_rd_addr; // @[Core.scala 34:23]
  wire [63:0] exereg_io_out_imm; // @[Core.scala 34:23]
  wire [63:0] exereg_io_out_op1; // @[Core.scala 34:23]
  wire [63:0] exereg_io_out_op2; // @[Core.scala 34:23]
  wire [6:0] exereg_io_out_fu_code; // @[Core.scala 34:23]
  wire [15:0] exereg_io_out_alu_code; // @[Core.scala 34:23]
  wire [7:0] exereg_io_out_bu_code; // @[Core.scala 34:23]
  wire [6:0] exereg_io_out_lu_code; // @[Core.scala 34:23]
  wire [3:0] exereg_io_out_su_code; // @[Core.scala 34:23]
  wire [1:0] exereg_io_out_mu_code; // @[Core.scala 34:23]
  wire [7:0] exereg_io_out_du_code; // @[Core.scala 34:23]
  wire [7:0] exereg_io_out_csru_code; // @[Core.scala 34:23]
  wire [4:0] exereg_io_out_rs1_addr; // @[Core.scala 34:23]
  wire  exereg_io_out_putch; // @[Core.scala 34:23]
  wire  memreg_clock; // @[Core.scala 35:23]
  wire  memreg_reset; // @[Core.scala 35:23]
  wire  memreg_io_en; // @[Core.scala 35:23]
  wire  memreg_io_in_valid; // @[Core.scala 35:23]
  wire [63:0] memreg_io_in_pc; // @[Core.scala 35:23]
  wire [31:0] memreg_io_in_inst; // @[Core.scala 35:23]
  wire  memreg_io_in_rd_en; // @[Core.scala 35:23]
  wire [4:0] memreg_io_in_rd_addr; // @[Core.scala 35:23]
  wire [63:0] memreg_io_in_imm; // @[Core.scala 35:23]
  wire [63:0] memreg_io_in_op1; // @[Core.scala 35:23]
  wire [63:0] memreg_io_in_op2; // @[Core.scala 35:23]
  wire [63:0] memreg_io_in_alu_out; // @[Core.scala 35:23]
  wire [63:0] memreg_io_in_bu_out; // @[Core.scala 35:23]
  wire [63:0] memreg_io_in_mu_out; // @[Core.scala 35:23]
  wire [63:0] memreg_io_in_du_out; // @[Core.scala 35:23]
  wire [63:0] memreg_io_in_csru_out; // @[Core.scala 35:23]
  wire [6:0] memreg_io_in_fu_code; // @[Core.scala 35:23]
  wire [6:0] memreg_io_in_lu_code; // @[Core.scala 35:23]
  wire [3:0] memreg_io_in_su_code; // @[Core.scala 35:23]
  wire  memreg_io_in_putch; // @[Core.scala 35:23]
  wire  memreg_io_in_csr_wen; // @[Core.scala 35:23]
  wire [11:0] memreg_io_in_csr_waddr; // @[Core.scala 35:23]
  wire [63:0] memreg_io_in_csr_wdata; // @[Core.scala 35:23]
  wire  memreg_io_out_valid; // @[Core.scala 35:23]
  wire [63:0] memreg_io_out_pc; // @[Core.scala 35:23]
  wire [31:0] memreg_io_out_inst; // @[Core.scala 35:23]
  wire  memreg_io_out_rd_en; // @[Core.scala 35:23]
  wire [4:0] memreg_io_out_rd_addr; // @[Core.scala 35:23]
  wire [63:0] memreg_io_out_imm; // @[Core.scala 35:23]
  wire [63:0] memreg_io_out_op1; // @[Core.scala 35:23]
  wire [63:0] memreg_io_out_op2; // @[Core.scala 35:23]
  wire [63:0] memreg_io_out_alu_out; // @[Core.scala 35:23]
  wire [63:0] memreg_io_out_bu_out; // @[Core.scala 35:23]
  wire [63:0] memreg_io_out_mu_out; // @[Core.scala 35:23]
  wire [63:0] memreg_io_out_du_out; // @[Core.scala 35:23]
  wire [63:0] memreg_io_out_csru_out; // @[Core.scala 35:23]
  wire [6:0] memreg_io_out_fu_code; // @[Core.scala 35:23]
  wire [6:0] memreg_io_out_lu_code; // @[Core.scala 35:23]
  wire [3:0] memreg_io_out_su_code; // @[Core.scala 35:23]
  wire  memreg_io_out_putch; // @[Core.scala 35:23]
  wire  memreg_io_out_csr_wen; // @[Core.scala 35:23]
  wire [11:0] memreg_io_out_csr_waddr; // @[Core.scala 35:23]
  wire [63:0] memreg_io_out_csr_wdata; // @[Core.scala 35:23]
  wire  wbreg_clock; // @[Core.scala 36:23]
  wire  wbreg_reset; // @[Core.scala 36:23]
  wire  wbreg_io_en; // @[Core.scala 36:23]
  wire  wbreg_io_in_valid; // @[Core.scala 36:23]
  wire [63:0] wbreg_io_in_pc; // @[Core.scala 36:23]
  wire [31:0] wbreg_io_in_inst; // @[Core.scala 36:23]
  wire  wbreg_io_in_rd_en; // @[Core.scala 36:23]
  wire [4:0] wbreg_io_in_rd_addr; // @[Core.scala 36:23]
  wire [63:0] wbreg_io_in_alu_out; // @[Core.scala 36:23]
  wire [63:0] wbreg_io_in_bu_out; // @[Core.scala 36:23]
  wire [63:0] wbreg_io_in_mu_out; // @[Core.scala 36:23]
  wire [63:0] wbreg_io_in_du_out; // @[Core.scala 36:23]
  wire [63:0] wbreg_io_in_csru_out; // @[Core.scala 36:23]
  wire [6:0] wbreg_io_in_fu_code; // @[Core.scala 36:23]
  wire [6:0] wbreg_io_in_lu_code; // @[Core.scala 36:23]
  wire [5:0] wbreg_io_in_lu_shift; // @[Core.scala 36:23]
  wire  wbreg_io_in_putch; // @[Core.scala 36:23]
  wire  wbreg_io_in_csr_wen; // @[Core.scala 36:23]
  wire [11:0] wbreg_io_in_csr_waddr; // @[Core.scala 36:23]
  wire [63:0] wbreg_io_in_csr_wdata; // @[Core.scala 36:23]
  wire  wbreg_io_in_csr_set_mtip; // @[Core.scala 36:23]
  wire  wbreg_io_in_csr_clear_mtip; // @[Core.scala 36:23]
  wire  wbreg_io_out_valid; // @[Core.scala 36:23]
  wire [63:0] wbreg_io_out_pc; // @[Core.scala 36:23]
  wire [31:0] wbreg_io_out_inst; // @[Core.scala 36:23]
  wire  wbreg_io_out_rd_en; // @[Core.scala 36:23]
  wire [4:0] wbreg_io_out_rd_addr; // @[Core.scala 36:23]
  wire [63:0] wbreg_io_out_alu_out; // @[Core.scala 36:23]
  wire [63:0] wbreg_io_out_bu_out; // @[Core.scala 36:23]
  wire [63:0] wbreg_io_out_mu_out; // @[Core.scala 36:23]
  wire [63:0] wbreg_io_out_du_out; // @[Core.scala 36:23]
  wire [63:0] wbreg_io_out_csru_out; // @[Core.scala 36:23]
  wire [6:0] wbreg_io_out_fu_code; // @[Core.scala 36:23]
  wire [6:0] wbreg_io_out_lu_code; // @[Core.scala 36:23]
  wire [5:0] wbreg_io_out_lu_shift; // @[Core.scala 36:23]
  wire  wbreg_io_out_putch; // @[Core.scala 36:23]
  wire  wbreg_io_out_csr_wen; // @[Core.scala 36:23]
  wire [11:0] wbreg_io_out_csr_waddr; // @[Core.scala 36:23]
  wire [63:0] wbreg_io_out_csr_wdata; // @[Core.scala 36:23]
  wire  wbreg_io_out_csr_set_mtip; // @[Core.scala 36:23]
  wire  wbreg_io_out_csr_clear_mtip; // @[Core.scala 36:23]
  wire  dt_ic_clock; // @[Core.scala 290:21]
  wire [7:0] dt_ic_coreid; // @[Core.scala 290:21]
  wire [7:0] dt_ic_index; // @[Core.scala 290:21]
  wire  dt_ic_valid; // @[Core.scala 290:21]
  wire [63:0] dt_ic_pc; // @[Core.scala 290:21]
  wire [31:0] dt_ic_instr; // @[Core.scala 290:21]
  wire [7:0] dt_ic_special; // @[Core.scala 290:21]
  wire  dt_ic_skip; // @[Core.scala 290:21]
  wire  dt_ic_isRVC; // @[Core.scala 290:21]
  wire  dt_ic_scFailed; // @[Core.scala 290:21]
  wire  dt_ic_wen; // @[Core.scala 290:21]
  wire [63:0] dt_ic_wdata; // @[Core.scala 290:21]
  wire [7:0] dt_ic_wdest; // @[Core.scala 290:21]
  wire  dt_ae_clock; // @[Core.scala 305:21]
  wire [7:0] dt_ae_coreid; // @[Core.scala 305:21]
  wire [31:0] dt_ae_intrNO; // @[Core.scala 305:21]
  wire [31:0] dt_ae_cause; // @[Core.scala 305:21]
  wire [63:0] dt_ae_exceptionPC; // @[Core.scala 305:21]
  wire [31:0] dt_ae_exceptionInst; // @[Core.scala 305:21]
  wire  dt_te_clock; // @[Core.scala 321:21]
  wire [7:0] dt_te_coreid; // @[Core.scala 321:21]
  wire  dt_te_valid; // @[Core.scala 321:21]
  wire [2:0] dt_te_code; // @[Core.scala 321:21]
  wire [63:0] dt_te_pc; // @[Core.scala 321:21]
  wire [63:0] dt_te_cycleCnt; // @[Core.scala 321:21]
  wire [63:0] dt_te_instrCnt; // @[Core.scala 321:21]
  wire  dmem_en = preamu_io_ren | preamu_io_wen; // @[Core.scala 126:31]
  wire  imem_not_ok = ~io_imem_ok; // @[Core.scala 209:21]
  wire  dmem_not_ok = ~io_dmem_ok; // @[Core.scala 210:21]
  wire [31:0] _exception_stall_T = idreg_io_inst; // @[Core.scala 215:40]
  wire  _exception_stall_T_1 = 32'h73 == _exception_stall_T; // @[Core.scala 215:40]
  wire  _exception_stall_T_3 = 32'h30200073 == _exception_stall_T; // @[Core.scala 215:67]
  wire  _exception_stall_T_4 = 32'h73 == _exception_stall_T | 32'h30200073 == _exception_stall_T; // @[Core.scala 215:50]
  wire  _exception_stall_T_6 = exereg_io_out_valid | memreg_io_out_valid | wbreg_io_out_valid; // @[Core.scala 215:124]
  wire  exception_stall = (32'h73 == _exception_stall_T | 32'h30200073 == _exception_stall_T) & (exereg_io_out_valid |
    memreg_io_out_valid | wbreg_io_out_valid); // @[Core.scala 215:77]
  wire  _fence_wait_T_1 = 32'h100f == _exception_stall_T; // @[Core.scala 226:34]
  wire  fence_wait = 32'h100f == _exception_stall_T & _exception_stall_T_6; // @[Core.scala 226:45]
  wire  fence_running = ~fence_io_ok; // @[Core.scala 228:23]
  wire  stall_id = rfconflict_io_conflict | imem_not_ok | exception_stall | fence_wait | fence_running; // @[Core.scala 238:86]
  wire  _exception_execution_T = ~stall_id; // @[Core.scala 216:29]
  wire  _exception_execution_T_7 = ~exereg_io_out_valid; // @[Core.scala 216:97]
  wire  _exception_execution_T_9 = ~memreg_io_out_valid; // @[Core.scala 216:121]
  wire  _exception_execution_T_11 = ~wbreg_io_out_valid; // @[Core.scala 216:145]
  wire  exception_execution = ~stall_id & _exception_stall_T_4 & ~exereg_io_out_valid & ~memreg_io_out_valid & ~
    wbreg_io_out_valid; // @[Core.scala 216:142]
  wire  stall_ie = mu_io_stall[0]; // @[Core.scala 207:22 Core.scala 241:12]
  wire  _memreg_io_in_valid_T = ~stall_ie; // @[Core.scala 251:48]
  wire  _commit_valid_T = ~dmem_not_ok; // @[Core.scala 253:44]
  wire  commit_valid = wbreg_io_out_valid & ~dmem_not_ok; // @[Core.scala 253:41]
  wire  skip_putch = wbreg_io_out_inst == 32'h7b; // @[Core.scala 278:38]
  wire [31:0] _read_mcycle_T = wbreg_io_out_inst & 32'hfff0307f; // @[Core.scala 279:27]
  wire  read_mcycle = _read_mcycle_T == 32'hb0002073; // @[Core.scala 279:44]
  wire  rtthread_test_skip = wbreg_io_out_inst == 32'h344737f3; // @[Core.scala 280:34]
  reg  skip_clint_REG; // @[Core.scala 281:35]
  reg  skip_clint; // @[Core.scala 281:27]
  reg  wbreg_exception_execution_REG; // @[Core.scala 284:66]
  reg  wbreg_exception_execution_REG_1; // @[Core.scala 284:58]
  reg  wbreg_exception_execution_REG_2; // @[Core.scala 284:50]
  reg  wbreg_exception_execution; // @[Core.scala 284:42]
  reg  wbreg_time_intr_REG; // @[Core.scala 285:66]
  reg  wbreg_time_intr_REG_1; // @[Core.scala 285:58]
  reg  wbreg_time_intr_REG_2; // @[Core.scala 285:50]
  reg  wbreg_time_intr; // @[Core.scala 285:42]
  reg [63:0] wbreg_cause_REG; // @[Core.scala 286:66]
  reg [63:0] wbreg_cause_REG_1; // @[Core.scala 286:58]
  reg [63:0] wbreg_cause_REG_2; // @[Core.scala 286:50]
  reg [63:0] wbreg_cause; // @[Core.scala 286:42]
  reg [63:0] wbreg_exception_pc_REG; // @[Core.scala 287:66]
  reg [63:0] wbreg_exception_pc_REG_1; // @[Core.scala 287:58]
  reg [63:0] wbreg_exception_pc_REG_2; // @[Core.scala 287:50]
  reg [63:0] wbreg_exception_pc; // @[Core.scala 287:42]
  wire [31:0] _commit_intr_T_1 = wbreg_io_out_inst; // @[Core.scala 288:82]
  reg  commit_intr_REG; // @[Core.scala 288:76]
  wire  commit_intr = wbreg_exception_execution & wbreg_time_intr & commit_intr_REG; // @[Core.scala 288:66]
  reg  dt_ic_io_valid_REG; // @[Core.scala 294:57]
  reg [63:0] dt_ic_io_pc_REG; // @[Core.scala 295:31]
  reg [31:0] dt_ic_io_instr_REG; // @[Core.scala 296:31]
  reg  dt_ic_io_skip_REG; // @[Core.scala 298:45]
  reg  dt_ic_io_wen_REG; // @[Core.scala 301:31]
  reg [63:0] dt_ic_io_wdata_REG; // @[Core.scala 302:31]
  reg [4:0] dt_ic_io_wdest_REG; // @[Core.scala 303:31]
  reg [63:0] cycle_cnt; // @[Core.scala 312:26]
  reg [63:0] instr_cnt; // @[Core.scala 313:26]
  wire [63:0] _cycle_cnt_T_1 = cycle_cnt + 64'h1; // @[Core.scala 315:26]
  wire [63:0] _instr_cnt_T_1 = instr_cnt + 64'h1; // @[Core.scala 316:44]
  wire [63:0] rf_a0_0 = rfu_rf_10;
  IFetch ifu ( // @[Core.scala 19:23]
    .reset(ifu_reset),
    .io_jump_en(ifu_io_jump_en),
    .io_jump_pc(ifu_io_jump_pc),
    .io_pc(ifu_io_pc),
    .io_next_pc(ifu_io_next_pc),
    .io_valid(ifu_io_valid)
  );
  Decode idu ( // @[Core.scala 20:23]
    .io_pc(idu_io_pc),
    .io_inst(idu_io_inst),
    .io_rs1_en(idu_io_rs1_en),
    .io_rs2_en(idu_io_rs2_en),
    .io_rs1_addr(idu_io_rs1_addr),
    .io_rs2_addr(idu_io_rs2_addr),
    .io_rs1_data(idu_io_rs1_data),
    .io_rs2_data(idu_io_rs2_data),
    .io_rd_en(idu_io_rd_en),
    .io_rd_addr(idu_io_rd_addr),
    .io_decode_info_fu_code(idu_io_decode_info_fu_code),
    .io_decode_info_alu_code(idu_io_decode_info_alu_code),
    .io_decode_info_bu_code(idu_io_decode_info_bu_code),
    .io_decode_info_lu_code(idu_io_decode_info_lu_code),
    .io_decode_info_su_code(idu_io_decode_info_su_code),
    .io_decode_info_mu_code(idu_io_decode_info_mu_code),
    .io_decode_info_du_code(idu_io_decode_info_du_code),
    .io_decode_info_csru_code(idu_io_decode_info_csru_code),
    .io_jump_en(idu_io_jump_en),
    .io_jump_pc(idu_io_jump_pc),
    .io_op1(idu_io_op1),
    .io_op2(idu_io_op2),
    .io_imm(idu_io_imm),
    .io_putch(idu_io_putch),
    .io_mtvec(idu_io_mtvec),
    .io_mepc(idu_io_mepc)
  );
  Execution ieu ( // @[Core.scala 21:23]
    .io_alu_code(ieu_io_alu_code),
    .io_bu_code(ieu_io_bu_code),
    .io_du_code(ieu_io_du_code),
    .io_csru_code(ieu_io_csru_code),
    .io_op1(ieu_io_op1),
    .io_op2(ieu_io_op2),
    .io_pc(ieu_io_pc),
    .io_alu_out(ieu_io_alu_out),
    .io_bu_out(ieu_io_bu_out),
    .io_du_out(ieu_io_du_out),
    .io_csru_out(ieu_io_csru_out),
    .io_rs1_addr(ieu_io_rs1_addr),
    .io_csr_raddr(ieu_io_csr_raddr),
    .io_csr_rdata(ieu_io_csr_rdata),
    .io_csr_wen(ieu_io_csr_wen),
    .io_csr_waddr(ieu_io_csr_waddr),
    .io_csr_wdata(ieu_io_csr_wdata)
  );
  RegFile rfu ( // @[Core.scala 22:23]
    .clock(rfu_clock),
    .reset(rfu_reset),
    .io_rs1_addr(rfu_io_rs1_addr),
    .io_rs2_addr(rfu_io_rs2_addr),
    .io_rs1_data(rfu_io_rs1_data),
    .io_rs2_data(rfu_io_rs2_data),
    .io_rd_addr(rfu_io_rd_addr),
    .io_rd_data(rfu_io_rd_data),
    .io_rd_en(rfu_io_rd_en),
    .rf_10(rfu_rf_10)
  );
  Csr csru ( // @[Core.scala 23:23]
    .clock(csru_clock),
    .reset(csru_reset),
    .io_raddr(csru_io_raddr),
    .io_rdata(csru_io_rdata),
    .io_wen(csru_io_wen),
    .io_waddr(csru_io_waddr),
    .io_wdata(csru_io_wdata),
    .io_set_mtip(csru_io_set_mtip),
    .io_clear_mtip(csru_io_clear_mtip),
    .io_exception(csru_io_exception),
    .io_cause(csru_io_cause),
    .io_mret(csru_io_mret),
    .io_pc(csru_io_pc),
    .io_mtvec(csru_io_mtvec),
    .io_mepc(csru_io_mepc),
    .io_time_intr(csru_io_time_intr)
  );
  PreAccessMemory preamu ( // @[Core.scala 24:23]
    .io_lu_code(preamu_io_lu_code),
    .io_su_code(preamu_io_su_code),
    .io_op1(preamu_io_op1),
    .io_op2(preamu_io_op2),
    .io_imm(preamu_io_imm),
    .io_lu_shift(preamu_io_lu_shift),
    .io_ren(preamu_io_ren),
    .io_raddr(preamu_io_raddr),
    .io_wen(preamu_io_wen),
    .io_waddr(preamu_io_waddr),
    .io_wdata(preamu_io_wdata),
    .io_wmask(preamu_io_wmask),
    .io_transfer(preamu_io_transfer)
  );
  AccessMemory amu ( // @[Core.scala 25:23]
    .io_lu_code(amu_io_lu_code),
    .io_lu_shift(amu_io_lu_shift),
    .io_rdata(amu_io_rdata),
    .io_lu_out(amu_io_lu_out)
  );
  WriteBack wbu ( // @[Core.scala 26:23]
    .io_fu_code(wbu_io_fu_code),
    .io_alu_out(wbu_io_alu_out),
    .io_bu_out(wbu_io_bu_out),
    .io_mu_out(wbu_io_mu_out),
    .io_du_out(wbu_io_du_out),
    .io_lu_out(wbu_io_lu_out),
    .io_csru_out(wbu_io_csru_out),
    .io_out(wbu_io_out)
  );
  MU mu ( // @[Core.scala 28:23]
    .clock(mu_clock),
    .reset(mu_reset),
    .io_en(mu_io_en),
    .io_mu_code(mu_io_mu_code),
    .io_op1(mu_io_op1),
    .io_op2(mu_io_op2),
    .io_mu_out(mu_io_mu_out),
    .io_stall(mu_io_stall)
  );
  RegfileConflict rfconflict ( // @[Core.scala 30:27]
    .io_rs_valid(rfconflict_io_rs_valid),
    .io_rs1_en(rfconflict_io_rs1_en),
    .io_rs2_en(rfconflict_io_rs2_en),
    .io_rs1_addr(rfconflict_io_rs1_addr),
    .io_rs2_addr(rfconflict_io_rs2_addr),
    .io_rd1_valid(rfconflict_io_rd1_valid),
    .io_rd1_en(rfconflict_io_rd1_en),
    .io_rd1_addr(rfconflict_io_rd1_addr),
    .io_rd2_valid(rfconflict_io_rd2_valid),
    .io_rd2_en(rfconflict_io_rd2_en),
    .io_rd2_addr(rfconflict_io_rd2_addr),
    .io_rd3_valid(rfconflict_io_rd3_valid),
    .io_rd3_en(rfconflict_io_rd3_en),
    .io_rd3_addr(rfconflict_io_rd3_addr),
    .io_conflict(rfconflict_io_conflict)
  );
  Fence fence ( // @[Core.scala 31:21]
    .clock(fence_clock),
    .reset(fence_reset),
    .io_go(fence_io_go),
    .io_ok(fence_io_ok),
    .io_ifence_req(fence_io_ifence_req),
    .io_ifence_done(fence_io_ifence_done),
    .io_dfence_req(fence_io_dfence_req),
    .io_dfence_done(fence_io_dfence_done)
  );
  IDReg idreg ( // @[Core.scala 33:23]
    .clock(idreg_clock),
    .reset(idreg_reset),
    .io_en(idreg_io_en),
    .io_in_valid(idreg_io_in_valid),
    .io_in_pc(idreg_io_in_pc),
    .io_out_valid(idreg_io_out_valid),
    .io_out_pc(idreg_io_out_pc),
    .io_imem__addr(idreg_io_imem__addr),
    .io_imem__en(idreg_io_imem__en),
    .io_imem__data(idreg_io_imem__data),
    .io_inst(idreg_io_inst)
  );
  ExeReg exereg ( // @[Core.scala 34:23]
    .clock(exereg_clock),
    .reset(exereg_reset),
    .io_en(exereg_io_en),
    .io_in_valid(exereg_io_in_valid),
    .io_in_pc(exereg_io_in_pc),
    .io_in_inst(exereg_io_in_inst),
    .io_in_rd_en(exereg_io_in_rd_en),
    .io_in_rd_addr(exereg_io_in_rd_addr),
    .io_in_imm(exereg_io_in_imm),
    .io_in_op1(exereg_io_in_op1),
    .io_in_op2(exereg_io_in_op2),
    .io_in_fu_code(exereg_io_in_fu_code),
    .io_in_alu_code(exereg_io_in_alu_code),
    .io_in_bu_code(exereg_io_in_bu_code),
    .io_in_lu_code(exereg_io_in_lu_code),
    .io_in_su_code(exereg_io_in_su_code),
    .io_in_mu_code(exereg_io_in_mu_code),
    .io_in_du_code(exereg_io_in_du_code),
    .io_in_csru_code(exereg_io_in_csru_code),
    .io_in_rs1_addr(exereg_io_in_rs1_addr),
    .io_in_putch(exereg_io_in_putch),
    .io_out_valid(exereg_io_out_valid),
    .io_out_pc(exereg_io_out_pc),
    .io_out_inst(exereg_io_out_inst),
    .io_out_rd_en(exereg_io_out_rd_en),
    .io_out_rd_addr(exereg_io_out_rd_addr),
    .io_out_imm(exereg_io_out_imm),
    .io_out_op1(exereg_io_out_op1),
    .io_out_op2(exereg_io_out_op2),
    .io_out_fu_code(exereg_io_out_fu_code),
    .io_out_alu_code(exereg_io_out_alu_code),
    .io_out_bu_code(exereg_io_out_bu_code),
    .io_out_lu_code(exereg_io_out_lu_code),
    .io_out_su_code(exereg_io_out_su_code),
    .io_out_mu_code(exereg_io_out_mu_code),
    .io_out_du_code(exereg_io_out_du_code),
    .io_out_csru_code(exereg_io_out_csru_code),
    .io_out_rs1_addr(exereg_io_out_rs1_addr),
    .io_out_putch(exereg_io_out_putch)
  );
  MemReg memreg ( // @[Core.scala 35:23]
    .clock(memreg_clock),
    .reset(memreg_reset),
    .io_en(memreg_io_en),
    .io_in_valid(memreg_io_in_valid),
    .io_in_pc(memreg_io_in_pc),
    .io_in_inst(memreg_io_in_inst),
    .io_in_rd_en(memreg_io_in_rd_en),
    .io_in_rd_addr(memreg_io_in_rd_addr),
    .io_in_imm(memreg_io_in_imm),
    .io_in_op1(memreg_io_in_op1),
    .io_in_op2(memreg_io_in_op2),
    .io_in_alu_out(memreg_io_in_alu_out),
    .io_in_bu_out(memreg_io_in_bu_out),
    .io_in_mu_out(memreg_io_in_mu_out),
    .io_in_du_out(memreg_io_in_du_out),
    .io_in_csru_out(memreg_io_in_csru_out),
    .io_in_fu_code(memreg_io_in_fu_code),
    .io_in_lu_code(memreg_io_in_lu_code),
    .io_in_su_code(memreg_io_in_su_code),
    .io_in_putch(memreg_io_in_putch),
    .io_in_csr_wen(memreg_io_in_csr_wen),
    .io_in_csr_waddr(memreg_io_in_csr_waddr),
    .io_in_csr_wdata(memreg_io_in_csr_wdata),
    .io_out_valid(memreg_io_out_valid),
    .io_out_pc(memreg_io_out_pc),
    .io_out_inst(memreg_io_out_inst),
    .io_out_rd_en(memreg_io_out_rd_en),
    .io_out_rd_addr(memreg_io_out_rd_addr),
    .io_out_imm(memreg_io_out_imm),
    .io_out_op1(memreg_io_out_op1),
    .io_out_op2(memreg_io_out_op2),
    .io_out_alu_out(memreg_io_out_alu_out),
    .io_out_bu_out(memreg_io_out_bu_out),
    .io_out_mu_out(memreg_io_out_mu_out),
    .io_out_du_out(memreg_io_out_du_out),
    .io_out_csru_out(memreg_io_out_csru_out),
    .io_out_fu_code(memreg_io_out_fu_code),
    .io_out_lu_code(memreg_io_out_lu_code),
    .io_out_su_code(memreg_io_out_su_code),
    .io_out_putch(memreg_io_out_putch),
    .io_out_csr_wen(memreg_io_out_csr_wen),
    .io_out_csr_waddr(memreg_io_out_csr_waddr),
    .io_out_csr_wdata(memreg_io_out_csr_wdata)
  );
  WBReg wbreg ( // @[Core.scala 36:23]
    .clock(wbreg_clock),
    .reset(wbreg_reset),
    .io_en(wbreg_io_en),
    .io_in_valid(wbreg_io_in_valid),
    .io_in_pc(wbreg_io_in_pc),
    .io_in_inst(wbreg_io_in_inst),
    .io_in_rd_en(wbreg_io_in_rd_en),
    .io_in_rd_addr(wbreg_io_in_rd_addr),
    .io_in_alu_out(wbreg_io_in_alu_out),
    .io_in_bu_out(wbreg_io_in_bu_out),
    .io_in_mu_out(wbreg_io_in_mu_out),
    .io_in_du_out(wbreg_io_in_du_out),
    .io_in_csru_out(wbreg_io_in_csru_out),
    .io_in_fu_code(wbreg_io_in_fu_code),
    .io_in_lu_code(wbreg_io_in_lu_code),
    .io_in_lu_shift(wbreg_io_in_lu_shift),
    .io_in_putch(wbreg_io_in_putch),
    .io_in_csr_wen(wbreg_io_in_csr_wen),
    .io_in_csr_waddr(wbreg_io_in_csr_waddr),
    .io_in_csr_wdata(wbreg_io_in_csr_wdata),
    .io_in_csr_set_mtip(wbreg_io_in_csr_set_mtip),
    .io_in_csr_clear_mtip(wbreg_io_in_csr_clear_mtip),
    .io_out_valid(wbreg_io_out_valid),
    .io_out_pc(wbreg_io_out_pc),
    .io_out_inst(wbreg_io_out_inst),
    .io_out_rd_en(wbreg_io_out_rd_en),
    .io_out_rd_addr(wbreg_io_out_rd_addr),
    .io_out_alu_out(wbreg_io_out_alu_out),
    .io_out_bu_out(wbreg_io_out_bu_out),
    .io_out_mu_out(wbreg_io_out_mu_out),
    .io_out_du_out(wbreg_io_out_du_out),
    .io_out_csru_out(wbreg_io_out_csru_out),
    .io_out_fu_code(wbreg_io_out_fu_code),
    .io_out_lu_code(wbreg_io_out_lu_code),
    .io_out_lu_shift(wbreg_io_out_lu_shift),
    .io_out_putch(wbreg_io_out_putch),
    .io_out_csr_wen(wbreg_io_out_csr_wen),
    .io_out_csr_waddr(wbreg_io_out_csr_waddr),
    .io_out_csr_wdata(wbreg_io_out_csr_wdata),
    .io_out_csr_set_mtip(wbreg_io_out_csr_set_mtip),
    .io_out_csr_clear_mtip(wbreg_io_out_csr_clear_mtip)
  );
  DifftestInstrCommit dt_ic ( // @[Core.scala 290:21]
    .clock(dt_ic_clock),
    .coreid(dt_ic_coreid),
    .index(dt_ic_index),
    .valid(dt_ic_valid),
    .pc(dt_ic_pc),
    .instr(dt_ic_instr),
    .special(dt_ic_special),
    .skip(dt_ic_skip),
    .isRVC(dt_ic_isRVC),
    .scFailed(dt_ic_scFailed),
    .wen(dt_ic_wen),
    .wdata(dt_ic_wdata),
    .wdest(dt_ic_wdest)
  );
  DifftestArchEvent dt_ae ( // @[Core.scala 305:21]
    .clock(dt_ae_clock),
    .coreid(dt_ae_coreid),
    .intrNO(dt_ae_intrNO),
    .cause(dt_ae_cause),
    .exceptionPC(dt_ae_exceptionPC),
    .exceptionInst(dt_ae_exceptionInst)
  );
  DifftestTrapEvent dt_te ( // @[Core.scala 321:21]
    .clock(dt_te_clock),
    .coreid(dt_te_coreid),
    .valid(dt_te_valid),
    .code(dt_te_code),
    .pc(dt_te_pc),
    .cycleCnt(dt_te_cycleCnt),
    .instrCnt(dt_te_instrCnt)
  );
  assign io_imem_addr = idreg_io_imem__addr; // @[Core.scala 42:17]
  assign io_imem_en = idreg_io_imem__en; // @[Core.scala 43:17]
  assign io_dmem_en = dmem_en & memreg_io_out_valid; // @[Core.scala 129:28]
  assign io_dmem_op = preamu_io_wen; // @[Core.scala 130:17]
  assign io_dmem_addr = preamu_io_wen ? preamu_io_waddr : preamu_io_raddr; // @[Core.scala 128:22]
  assign io_dmem_wdata = preamu_io_wdata; // @[Core.scala 132:17]
  assign io_dmem_wmask = preamu_io_wmask; // @[Core.scala 133:17]
  assign io_dmem_transfer = {{29'd0}, preamu_io_transfer}; // @[Core.scala 134:20]
  assign io_ifence_req = fence_io_ifence_req; // @[Core.scala 230:19]
  assign io_dfence_req = fence_io_dfence_req; // @[Core.scala 231:19]
  assign ifu_reset = reset;
  assign ifu_io_jump_en = idu_io_jump_en; // @[Core.scala 38:19]
  assign ifu_io_jump_pc = idu_io_jump_pc; // @[Core.scala 39:19]
  assign ifu_io_pc = idreg_io_out_pc; // @[Core.scala 40:19]
  assign idu_io_pc = idreg_io_out_pc; // @[Core.scala 49:19]
  assign idu_io_inst = idreg_io_inst; // @[Core.scala 50:19]
  assign idu_io_rs1_data = rfu_io_rs1_data; // @[Core.scala 51:19]
  assign idu_io_rs2_data = rfu_io_rs2_data; // @[Core.scala 52:19]
  assign idu_io_mtvec = csru_io_mtvec; // @[Core.scala 53:19]
  assign idu_io_mepc = csru_io_mepc; // @[Core.scala 54:19]
  assign ieu_io_alu_code = exereg_io_out_alu_code; // @[Core.scala 75:21]
  assign ieu_io_bu_code = exereg_io_out_bu_code; // @[Core.scala 76:21]
  assign ieu_io_du_code = exereg_io_out_du_code; // @[Core.scala 77:21]
  assign ieu_io_csru_code = exereg_io_out_csru_code; // @[Core.scala 80:21]
  assign ieu_io_op1 = exereg_io_out_op1; // @[Core.scala 81:14]
  assign ieu_io_op2 = exereg_io_out_op2; // @[Core.scala 82:14]
  assign ieu_io_pc = exereg_io_out_pc; // @[Core.scala 83:14]
  assign ieu_io_rs1_addr = exereg_io_out_rs1_addr; // @[Core.scala 85:19]
  assign ieu_io_csr_rdata = csru_io_rdata; // @[Core.scala 86:20]
  assign rfu_clock = clock;
  assign rfu_reset = reset;
  assign rfu_io_rs1_addr = idu_io_rs1_addr; // @[Core.scala 174:19]
  assign rfu_io_rs2_addr = idu_io_rs2_addr; // @[Core.scala 175:19]
  assign rfu_io_rd_addr = wbreg_io_out_rd_addr; // @[Core.scala 177:19]
  assign rfu_io_rd_data = wbu_io_out; // @[Core.scala 179:19]
  assign rfu_io_rd_en = wbreg_io_out_rd_en & commit_valid; // @[Core.scala 261:39]
  assign csru_clock = clock;
  assign csru_reset = reset;
  assign csru_io_raddr = ieu_io_csr_raddr; // @[Core.scala 182:21]
  assign csru_io_wen = wbreg_io_out_csr_wen & commit_valid; // @[Core.scala 262:41]
  assign csru_io_waddr = wbreg_io_out_csr_waddr; // @[Core.scala 183:21]
  assign csru_io_wdata = wbreg_io_out_csr_wdata; // @[Core.scala 184:21]
  assign csru_io_set_mtip = wbreg_io_out_csr_set_mtip; // @[Core.scala 186:23]
  assign csru_io_clear_mtip = wbreg_io_out_csr_clear_mtip; // @[Core.scala 187:23]
  assign csru_io_exception = exception_execution & _exception_stall_T_1; // @[Core.scala 217:44]
  assign csru_io_cause = csru_io_time_intr ? 64'h8000000000000007 : 64'hb; // @[Core.scala 219:27]
  assign csru_io_mret = exception_execution & _exception_stall_T_3; // @[Core.scala 218:44]
  assign csru_io_pc = idreg_io_out_pc; // @[Core.scala 220:21]
  assign preamu_io_lu_code = memreg_io_out_lu_code; // @[Core.scala 120:21]
  assign preamu_io_su_code = memreg_io_out_su_code; // @[Core.scala 121:21]
  assign preamu_io_op1 = memreg_io_out_op1; // @[Core.scala 122:21]
  assign preamu_io_op2 = memreg_io_out_op2; // @[Core.scala 123:21]
  assign preamu_io_imm = memreg_io_out_imm; // @[Core.scala 124:21]
  assign amu_io_lu_code = wbreg_io_out_lu_code; // @[Core.scala 159:19]
  assign amu_io_lu_shift = wbreg_io_out_lu_shift; // @[Core.scala 160:19]
  assign amu_io_rdata = io_dmem_rdata; // @[Core.scala 161:19]
  assign wbu_io_fu_code = wbreg_io_out_fu_code; // @[Core.scala 163:19]
  assign wbu_io_alu_out = wbreg_io_out_alu_out; // @[Core.scala 164:19]
  assign wbu_io_bu_out = wbreg_io_out_bu_out; // @[Core.scala 165:19]
  assign wbu_io_mu_out = wbreg_io_out_mu_out; // @[Core.scala 166:19]
  assign wbu_io_du_out = wbreg_io_out_du_out; // @[Core.scala 167:19]
  assign wbu_io_lu_out = amu_io_lu_out; // @[Core.scala 169:19]
  assign wbu_io_csru_out = wbreg_io_out_csru_out; // @[Core.scala 168:19]
  assign mu_clock = clock;
  assign mu_reset = reset;
  assign mu_io_en = exereg_io_out_valid & exereg_io_out_mu_code != 2'h0; // @[Core.scala 88:40]
  assign mu_io_mu_code = exereg_io_out_mu_code; // @[Core.scala 89:17]
  assign mu_io_op1 = exereg_io_out_op1; // @[Core.scala 90:17]
  assign mu_io_op2 = exereg_io_out_op2; // @[Core.scala 91:17]
  assign rfconflict_io_rs_valid = idreg_io_out_valid; // @[Core.scala 190:28]
  assign rfconflict_io_rs1_en = idu_io_rs1_en; // @[Core.scala 191:28]
  assign rfconflict_io_rs2_en = idu_io_rs2_en; // @[Core.scala 192:28]
  assign rfconflict_io_rs1_addr = idu_io_rs1_addr; // @[Core.scala 193:28]
  assign rfconflict_io_rs2_addr = idu_io_rs2_addr; // @[Core.scala 194:28]
  assign rfconflict_io_rd1_valid = exereg_io_out_valid; // @[Core.scala 195:28]
  assign rfconflict_io_rd1_en = exereg_io_out_rd_en; // @[Core.scala 196:28]
  assign rfconflict_io_rd1_addr = exereg_io_out_rd_addr; // @[Core.scala 197:28]
  assign rfconflict_io_rd2_valid = memreg_io_out_valid; // @[Core.scala 198:28]
  assign rfconflict_io_rd2_en = memreg_io_out_rd_en; // @[Core.scala 199:28]
  assign rfconflict_io_rd2_addr = memreg_io_out_rd_addr; // @[Core.scala 200:28]
  assign rfconflict_io_rd3_valid = wbreg_io_out_valid; // @[Core.scala 201:28]
  assign rfconflict_io_rd3_en = wbreg_io_out_rd_en; // @[Core.scala 202:28]
  assign rfconflict_io_rd3_addr = wbreg_io_out_rd_addr; // @[Core.scala 203:28]
  assign fence_clock = clock;
  assign fence_reset = reset;
  assign fence_io_go = _fence_wait_T_1 & _exception_execution_T_7 & _exception_execution_T_9 & _exception_execution_T_11
    ; // @[Core.scala 227:91]
  assign fence_io_ifence_done = io_ifence_done; // @[Core.scala 230:19]
  assign fence_io_dfence_done = io_dfence_done; // @[Core.scala 231:19]
  assign idreg_clock = clock;
  assign idreg_reset = reset;
  assign idreg_io_en = _commit_valid_T & _memreg_io_in_valid_T & _exception_execution_T; // @[Core.scala 255:42]
  assign idreg_io_in_valid = ifu_io_valid; // @[Core.scala 249:22]
  assign idreg_io_in_pc = ifu_io_next_pc; // @[Core.scala 47:19]
  assign idreg_io_imem__data = csru_io_time_intr ? 32'h73 : io_imem_data; // @[Core.scala 222:29]
  assign exereg_clock = clock;
  assign exereg_reset = reset;
  assign exereg_io_en = _commit_valid_T & _memreg_io_in_valid_T; // @[Core.scala 256:29]
  assign exereg_io_in_valid = idreg_io_out_valid & _exception_execution_T; // @[Core.scala 250:44]
  assign exereg_io_in_pc = idreg_io_out_pc; // @[Core.scala 56:27]
  assign exereg_io_in_inst = idreg_io_inst; // @[Core.scala 57:27]
  assign exereg_io_in_rd_en = idu_io_rd_en; // @[Core.scala 58:27]
  assign exereg_io_in_rd_addr = idu_io_rd_addr; // @[Core.scala 59:27]
  assign exereg_io_in_imm = idu_io_imm; // @[Core.scala 60:27]
  assign exereg_io_in_op1 = idu_io_op1; // @[Core.scala 61:27]
  assign exereg_io_in_op2 = idu_io_op2; // @[Core.scala 62:27]
  assign exereg_io_in_fu_code = idu_io_decode_info_fu_code; // @[Core.scala 64:27]
  assign exereg_io_in_alu_code = idu_io_decode_info_alu_code; // @[Core.scala 65:27]
  assign exereg_io_in_bu_code = idu_io_decode_info_bu_code; // @[Core.scala 66:27]
  assign exereg_io_in_lu_code = idu_io_decode_info_lu_code; // @[Core.scala 69:27]
  assign exereg_io_in_su_code = idu_io_decode_info_su_code; // @[Core.scala 70:27]
  assign exereg_io_in_mu_code = idu_io_decode_info_mu_code; // @[Core.scala 67:27]
  assign exereg_io_in_du_code = idu_io_decode_info_du_code; // @[Core.scala 68:27]
  assign exereg_io_in_csru_code = idu_io_decode_info_csru_code; // @[Core.scala 71:27]
  assign exereg_io_in_rs1_addr = idu_io_rs1_addr; // @[Core.scala 63:27]
  assign exereg_io_in_putch = idu_io_putch; // @[Core.scala 72:27]
  assign memreg_clock = clock;
  assign memreg_reset = reset;
  assign memreg_io_en = ~dmem_not_ok; // @[Core.scala 257:19]
  assign memreg_io_in_valid = exereg_io_out_valid & ~stall_ie; // @[Core.scala 251:45]
  assign memreg_io_in_pc = exereg_io_out_pc; // @[Core.scala 93:25]
  assign memreg_io_in_inst = exereg_io_out_inst; // @[Core.scala 94:25]
  assign memreg_io_in_rd_en = exereg_io_out_rd_en; // @[Core.scala 95:25]
  assign memreg_io_in_rd_addr = exereg_io_out_rd_addr; // @[Core.scala 96:25]
  assign memreg_io_in_imm = exereg_io_out_imm; // @[Core.scala 97:25]
  assign memreg_io_in_op1 = exereg_io_out_op1; // @[Core.scala 98:25]
  assign memreg_io_in_op2 = exereg_io_out_op2; // @[Core.scala 99:25]
  assign memreg_io_in_alu_out = ieu_io_alu_out; // @[Core.scala 109:25]
  assign memreg_io_in_bu_out = ieu_io_bu_out; // @[Core.scala 110:25]
  assign memreg_io_in_mu_out = mu_io_mu_out; // @[Core.scala 111:25]
  assign memreg_io_in_du_out = ieu_io_du_out; // @[Core.scala 112:25]
  assign memreg_io_in_csru_out = ieu_io_csru_out; // @[Core.scala 113:25]
  assign memreg_io_in_fu_code = exereg_io_out_fu_code; // @[Core.scala 100:25]
  assign memreg_io_in_lu_code = exereg_io_out_lu_code; // @[Core.scala 105:25]
  assign memreg_io_in_su_code = exereg_io_out_su_code; // @[Core.scala 106:25]
  assign memreg_io_in_putch = exereg_io_out_putch; // @[Core.scala 115:27]
  assign memreg_io_in_csr_wen = ieu_io_csr_wen; // @[Core.scala 116:27]
  assign memreg_io_in_csr_waddr = ieu_io_csr_waddr; // @[Core.scala 117:27]
  assign memreg_io_in_csr_wdata = ieu_io_csr_wdata; // @[Core.scala 118:27]
  assign wbreg_clock = clock;
  assign wbreg_reset = reset;
  assign wbreg_io_en = ~dmem_not_ok; // @[Core.scala 258:19]
  assign wbreg_io_in_valid = memreg_io_out_valid; // @[Core.scala 252:22]
  assign wbreg_io_in_pc = memreg_io_out_pc; // @[Core.scala 136:25]
  assign wbreg_io_in_inst = memreg_io_out_inst; // @[Core.scala 137:25]
  assign wbreg_io_in_rd_en = memreg_io_out_rd_en; // @[Core.scala 138:25]
  assign wbreg_io_in_rd_addr = memreg_io_out_rd_addr; // @[Core.scala 139:25]
  assign wbreg_io_in_alu_out = memreg_io_out_alu_out; // @[Core.scala 140:25]
  assign wbreg_io_in_bu_out = memreg_io_out_bu_out; // @[Core.scala 141:25]
  assign wbreg_io_in_mu_out = memreg_io_out_mu_out; // @[Core.scala 142:25]
  assign wbreg_io_in_du_out = memreg_io_out_du_out; // @[Core.scala 143:25]
  assign wbreg_io_in_csru_out = memreg_io_out_csru_out; // @[Core.scala 144:25]
  assign wbreg_io_in_fu_code = memreg_io_out_fu_code; // @[Core.scala 145:25]
  assign wbreg_io_in_lu_code = memreg_io_out_lu_code; // @[Core.scala 146:25]
  assign wbreg_io_in_lu_shift = preamu_io_lu_shift; // @[Core.scala 149:25]
  assign wbreg_io_in_putch = memreg_io_out_putch; // @[Core.scala 151:25]
  assign wbreg_io_in_csr_wen = memreg_io_out_csr_wen; // @[Core.scala 152:25]
  assign wbreg_io_in_csr_waddr = memreg_io_out_csr_waddr; // @[Core.scala 153:25]
  assign wbreg_io_in_csr_wdata = memreg_io_out_csr_wdata; // @[Core.scala 154:25]
  assign wbreg_io_in_csr_set_mtip = io_set_mtip; // @[Core.scala 156:31]
  assign wbreg_io_in_csr_clear_mtip = io_clear_mtip; // @[Core.scala 157:31]
  assign dt_ic_clock = clock; // @[Core.scala 291:21]
  assign dt_ic_coreid = 8'h0; // @[Core.scala 292:21]
  assign dt_ic_index = 8'h0; // @[Core.scala 293:21]
  assign dt_ic_valid = commit_intr ? 1'h0 : dt_ic_io_valid_REG; // @[Core.scala 294:27]
  assign dt_ic_pc = dt_ic_io_pc_REG; // @[Core.scala 295:21]
  assign dt_ic_instr = dt_ic_io_instr_REG; // @[Core.scala 296:21]
  assign dt_ic_special = 8'h0; // @[Core.scala 297:21]
  assign dt_ic_skip = skip_clint | dt_ic_io_skip_REG; // @[Core.scala 298:35]
  assign dt_ic_isRVC = 1'h0; // @[Core.scala 299:21]
  assign dt_ic_scFailed = 1'h0; // @[Core.scala 300:21]
  assign dt_ic_wen = dt_ic_io_wen_REG; // @[Core.scala 301:21]
  assign dt_ic_wdata = dt_ic_io_wdata_REG; // @[Core.scala 302:21]
  assign dt_ic_wdest = {{3'd0}, dt_ic_io_wdest_REG}; // @[Core.scala 303:21]
  assign dt_ae_clock = clock; // @[Core.scala 306:25]
  assign dt_ae_coreid = 8'h0; // @[Core.scala 307:25]
  assign dt_ae_intrNO = commit_intr ? wbreg_cause[31:0] : 32'h0; // @[Core.scala 308:31]
  assign dt_ae_cause = commit_intr ? wbreg_cause[31:0] : 32'h0; // @[Core.scala 309:31]
  assign dt_ae_exceptionPC = commit_intr ? wbreg_exception_pc : 64'h0; // @[Core.scala 310:31]
  assign dt_ae_exceptionInst = 32'h0;
  assign dt_te_clock = clock; // @[Core.scala 322:21]
  assign dt_te_coreid = 8'h0; // @[Core.scala 323:21]
  assign dt_te_valid = (wbreg_io_out_inst == 32'h6b | wbreg_io_out_inst == 32'h100073) & commit_valid; // @[Core.scala 324:101]
  assign dt_te_code = rf_a0_0[2:0]; // @[Core.scala 325:29]
  assign dt_te_pc = wbreg_io_out_pc; // @[Core.scala 326:21]
  assign dt_te_cycleCnt = cycle_cnt; // @[Core.scala 327:21]
  assign dt_te_instrCnt = instr_cnt; // @[Core.scala 328:21]
  always @(posedge clock) begin
    skip_clint_REG <= io_dmem_en & (io_dmem_addr == 64'h200bff8 | io_dmem_addr == 64'h2004000); // @[Core.scala 281:47]
    skip_clint <= skip_clint_REG; // @[Core.scala 281:27]
    wbreg_exception_execution_REG <= ~stall_id & _exception_stall_T_4 & ~exereg_io_out_valid & ~memreg_io_out_valid & ~
      wbreg_io_out_valid; // @[Core.scala 216:142]
    wbreg_exception_execution_REG_1 <= wbreg_exception_execution_REG; // @[Core.scala 284:58]
    wbreg_exception_execution_REG_2 <= wbreg_exception_execution_REG_1; // @[Core.scala 284:50]
    wbreg_exception_execution <= wbreg_exception_execution_REG_2; // @[Core.scala 284:42]
    wbreg_time_intr_REG <= csru_io_time_intr; // @[Core.scala 285:66]
    wbreg_time_intr_REG_1 <= wbreg_time_intr_REG; // @[Core.scala 285:58]
    wbreg_time_intr_REG_2 <= wbreg_time_intr_REG_1; // @[Core.scala 285:50]
    wbreg_time_intr <= wbreg_time_intr_REG_2; // @[Core.scala 285:42]
    wbreg_cause_REG <= csru_io_cause; // @[Core.scala 286:66]
    wbreg_cause_REG_1 <= wbreg_cause_REG; // @[Core.scala 286:58]
    wbreg_cause_REG_2 <= wbreg_cause_REG_1; // @[Core.scala 286:50]
    wbreg_cause <= wbreg_cause_REG_2; // @[Core.scala 286:42]
    wbreg_exception_pc_REG <= csru_io_pc; // @[Core.scala 287:66]
    wbreg_exception_pc_REG_1 <= wbreg_exception_pc_REG; // @[Core.scala 287:58]
    wbreg_exception_pc_REG_2 <= wbreg_exception_pc_REG_1; // @[Core.scala 287:50]
    wbreg_exception_pc <= wbreg_exception_pc_REG_2; // @[Core.scala 287:42]
    commit_intr_REG <= 32'h73 == _commit_intr_T_1; // @[Core.scala 288:82]
    dt_ic_io_valid_REG <= wbreg_io_out_valid & ~dmem_not_ok; // @[Core.scala 253:41]
    dt_ic_io_pc_REG <= wbreg_io_out_pc; // @[Core.scala 295:31]
    dt_ic_io_instr_REG <= wbreg_io_out_inst; // @[Core.scala 296:31]
    dt_ic_io_skip_REG <= skip_putch | read_mcycle | rtthread_test_skip; // @[Core.scala 298:72]
    dt_ic_io_wen_REG <= wbreg_io_out_rd_en; // @[Core.scala 301:31]
    dt_ic_io_wdata_REG <= wbu_io_out; // @[Core.scala 302:31]
    dt_ic_io_wdest_REG <= wbreg_io_out_rd_addr; // @[Core.scala 303:31]
    if (reset) begin // @[Core.scala 312:26]
      cycle_cnt <= 64'h0; // @[Core.scala 312:26]
    end else begin
      cycle_cnt <= _cycle_cnt_T_1; // @[Core.scala 315:13]
    end
    if (reset) begin // @[Core.scala 313:26]
      instr_cnt <= 64'h0; // @[Core.scala 313:26]
    end else if (commit_valid) begin // @[Core.scala 316:19]
      instr_cnt <= _instr_cnt_T_1;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (wbreg_io_out_putch & commit_valid & ~reset) begin
          $fwrite(32'h80000002,"%c",rf_a0_0); // @[Core.scala 271:51]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  skip_clint_REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  skip_clint = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  wbreg_exception_execution_REG = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  wbreg_exception_execution_REG_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  wbreg_exception_execution_REG_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  wbreg_exception_execution = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  wbreg_time_intr_REG = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  wbreg_time_intr_REG_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  wbreg_time_intr_REG_2 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  wbreg_time_intr = _RAND_9[0:0];
  _RAND_10 = {2{`RANDOM}};
  wbreg_cause_REG = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  wbreg_cause_REG_1 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  wbreg_cause_REG_2 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  wbreg_cause = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  wbreg_exception_pc_REG = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  wbreg_exception_pc_REG_1 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  wbreg_exception_pc_REG_2 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  wbreg_exception_pc = _RAND_17[63:0];
  _RAND_18 = {1{`RANDOM}};
  commit_intr_REG = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  dt_ic_io_valid_REG = _RAND_19[0:0];
  _RAND_20 = {2{`RANDOM}};
  dt_ic_io_pc_REG = _RAND_20[63:0];
  _RAND_21 = {1{`RANDOM}};
  dt_ic_io_instr_REG = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  dt_ic_io_skip_REG = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  dt_ic_io_wen_REG = _RAND_23[0:0];
  _RAND_24 = {2{`RANDOM}};
  dt_ic_io_wdata_REG = _RAND_24[63:0];
  _RAND_25 = {1{`RANDOM}};
  dt_ic_io_wdest_REG = _RAND_25[4:0];
  _RAND_26 = {2{`RANDOM}};
  cycle_cnt = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  instr_cnt = _RAND_27[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ICache(
  input          clock,
  input          reset,
  input  [63:0]  io_imem_addr,
  input          io_imem_en,
  output [31:0]  io_imem_data,
  output         io_imem_ok,
  output         io_axi_req,
  output [63:0]  io_axi_addr,
  input          io_axi_valid,
  input  [511:0] io_axi_data,
  input          io_fence_req,
  output         io_fence_done
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [63:0] _RAND_65;
  reg [63:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [63:0] _RAND_68;
  reg [63:0] _RAND_69;
  reg [63:0] _RAND_70;
  reg [63:0] _RAND_71;
  reg [63:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [63:0] _RAND_75;
  reg [63:0] _RAND_76;
  reg [63:0] _RAND_77;
  reg [63:0] _RAND_78;
  reg [63:0] _RAND_79;
  reg [63:0] _RAND_80;
  reg [63:0] _RAND_81;
  reg [63:0] _RAND_82;
  reg [63:0] _RAND_83;
  reg [63:0] _RAND_84;
  reg [63:0] _RAND_85;
  reg [63:0] _RAND_86;
  reg [63:0] _RAND_87;
  reg [63:0] _RAND_88;
  reg [63:0] _RAND_89;
  reg [63:0] _RAND_90;
  reg [63:0] _RAND_91;
  reg [63:0] _RAND_92;
  reg [63:0] _RAND_93;
  reg [63:0] _RAND_94;
  reg [63:0] _RAND_95;
  reg [63:0] _RAND_96;
  reg [511:0] _RAND_97;
  reg [511:0] _RAND_98;
  reg [511:0] _RAND_99;
  reg [511:0] _RAND_100;
  reg [511:0] _RAND_101;
  reg [511:0] _RAND_102;
  reg [511:0] _RAND_103;
  reg [511:0] _RAND_104;
  reg [511:0] _RAND_105;
  reg [511:0] _RAND_106;
  reg [511:0] _RAND_107;
  reg [511:0] _RAND_108;
  reg [511:0] _RAND_109;
  reg [511:0] _RAND_110;
  reg [511:0] _RAND_111;
  reg [511:0] _RAND_112;
  reg [511:0] _RAND_113;
  reg [511:0] _RAND_114;
  reg [511:0] _RAND_115;
  reg [511:0] _RAND_116;
  reg [511:0] _RAND_117;
  reg [511:0] _RAND_118;
  reg [511:0] _RAND_119;
  reg [511:0] _RAND_120;
  reg [511:0] _RAND_121;
  reg [511:0] _RAND_122;
  reg [511:0] _RAND_123;
  reg [511:0] _RAND_124;
  reg [511:0] _RAND_125;
  reg [511:0] _RAND_126;
  reg [511:0] _RAND_127;
  reg [511:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [63:0] _RAND_193;
  reg [63:0] _RAND_194;
  reg [63:0] _RAND_195;
  reg [63:0] _RAND_196;
  reg [63:0] _RAND_197;
  reg [63:0] _RAND_198;
  reg [63:0] _RAND_199;
  reg [63:0] _RAND_200;
  reg [63:0] _RAND_201;
  reg [63:0] _RAND_202;
  reg [63:0] _RAND_203;
  reg [63:0] _RAND_204;
  reg [63:0] _RAND_205;
  reg [63:0] _RAND_206;
  reg [63:0] _RAND_207;
  reg [63:0] _RAND_208;
  reg [63:0] _RAND_209;
  reg [63:0] _RAND_210;
  reg [63:0] _RAND_211;
  reg [63:0] _RAND_212;
  reg [63:0] _RAND_213;
  reg [63:0] _RAND_214;
  reg [63:0] _RAND_215;
  reg [63:0] _RAND_216;
  reg [63:0] _RAND_217;
  reg [63:0] _RAND_218;
  reg [63:0] _RAND_219;
  reg [63:0] _RAND_220;
  reg [63:0] _RAND_221;
  reg [63:0] _RAND_222;
  reg [63:0] _RAND_223;
  reg [63:0] _RAND_224;
  reg [511:0] _RAND_225;
  reg [511:0] _RAND_226;
  reg [511:0] _RAND_227;
  reg [511:0] _RAND_228;
  reg [511:0] _RAND_229;
  reg [511:0] _RAND_230;
  reg [511:0] _RAND_231;
  reg [511:0] _RAND_232;
  reg [511:0] _RAND_233;
  reg [511:0] _RAND_234;
  reg [511:0] _RAND_235;
  reg [511:0] _RAND_236;
  reg [511:0] _RAND_237;
  reg [511:0] _RAND_238;
  reg [511:0] _RAND_239;
  reg [511:0] _RAND_240;
  reg [511:0] _RAND_241;
  reg [511:0] _RAND_242;
  reg [511:0] _RAND_243;
  reg [511:0] _RAND_244;
  reg [511:0] _RAND_245;
  reg [511:0] _RAND_246;
  reg [511:0] _RAND_247;
  reg [511:0] _RAND_248;
  reg [511:0] _RAND_249;
  reg [511:0] _RAND_250;
  reg [511:0] _RAND_251;
  reg [511:0] _RAND_252;
  reg [511:0] _RAND_253;
  reg [511:0] _RAND_254;
  reg [511:0] _RAND_255;
  reg [511:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
`endif // RANDOMIZE_REG_INIT
  wire  _addr_T = io_imem_en & io_imem_ok; // @[ICache.scala 46:62]
  reg [63:0] addr; // @[Reg.scala 27:20]
  wire [52:0] tag_addr = addr[63:11]; // @[ICache.scala 49:27]
  wire [4:0] index_addr = addr[10:6]; // @[ICache.scala 50:27]
  wire [5:0] offset_addr = addr[5:0]; // @[ICache.scala 51:27]
  reg  v1_0; // @[ICache.scala 53:26]
  reg  v1_1; // @[ICache.scala 53:26]
  reg  v1_2; // @[ICache.scala 53:26]
  reg  v1_3; // @[ICache.scala 53:26]
  reg  v1_4; // @[ICache.scala 53:26]
  reg  v1_5; // @[ICache.scala 53:26]
  reg  v1_6; // @[ICache.scala 53:26]
  reg  v1_7; // @[ICache.scala 53:26]
  reg  v1_8; // @[ICache.scala 53:26]
  reg  v1_9; // @[ICache.scala 53:26]
  reg  v1_10; // @[ICache.scala 53:26]
  reg  v1_11; // @[ICache.scala 53:26]
  reg  v1_12; // @[ICache.scala 53:26]
  reg  v1_13; // @[ICache.scala 53:26]
  reg  v1_14; // @[ICache.scala 53:26]
  reg  v1_15; // @[ICache.scala 53:26]
  reg  v1_16; // @[ICache.scala 53:26]
  reg  v1_17; // @[ICache.scala 53:26]
  reg  v1_18; // @[ICache.scala 53:26]
  reg  v1_19; // @[ICache.scala 53:26]
  reg  v1_20; // @[ICache.scala 53:26]
  reg  v1_21; // @[ICache.scala 53:26]
  reg  v1_22; // @[ICache.scala 53:26]
  reg  v1_23; // @[ICache.scala 53:26]
  reg  v1_24; // @[ICache.scala 53:26]
  reg  v1_25; // @[ICache.scala 53:26]
  reg  v1_26; // @[ICache.scala 53:26]
  reg  v1_27; // @[ICache.scala 53:26]
  reg  v1_28; // @[ICache.scala 53:26]
  reg  v1_29; // @[ICache.scala 53:26]
  reg  v1_30; // @[ICache.scala 53:26]
  reg  v1_31; // @[ICache.scala 53:26]
  reg  age1_0; // @[ICache.scala 54:26]
  reg  age1_1; // @[ICache.scala 54:26]
  reg  age1_2; // @[ICache.scala 54:26]
  reg  age1_3; // @[ICache.scala 54:26]
  reg  age1_4; // @[ICache.scala 54:26]
  reg  age1_5; // @[ICache.scala 54:26]
  reg  age1_6; // @[ICache.scala 54:26]
  reg  age1_7; // @[ICache.scala 54:26]
  reg  age1_8; // @[ICache.scala 54:26]
  reg  age1_9; // @[ICache.scala 54:26]
  reg  age1_10; // @[ICache.scala 54:26]
  reg  age1_11; // @[ICache.scala 54:26]
  reg  age1_12; // @[ICache.scala 54:26]
  reg  age1_13; // @[ICache.scala 54:26]
  reg  age1_14; // @[ICache.scala 54:26]
  reg  age1_15; // @[ICache.scala 54:26]
  reg  age1_16; // @[ICache.scala 54:26]
  reg  age1_17; // @[ICache.scala 54:26]
  reg  age1_18; // @[ICache.scala 54:26]
  reg  age1_19; // @[ICache.scala 54:26]
  reg  age1_20; // @[ICache.scala 54:26]
  reg  age1_21; // @[ICache.scala 54:26]
  reg  age1_22; // @[ICache.scala 54:26]
  reg  age1_23; // @[ICache.scala 54:26]
  reg  age1_24; // @[ICache.scala 54:26]
  reg  age1_25; // @[ICache.scala 54:26]
  reg  age1_26; // @[ICache.scala 54:26]
  reg  age1_27; // @[ICache.scala 54:26]
  reg  age1_28; // @[ICache.scala 54:26]
  reg  age1_29; // @[ICache.scala 54:26]
  reg  age1_30; // @[ICache.scala 54:26]
  reg  age1_31; // @[ICache.scala 54:26]
  reg [52:0] tag1_0; // @[ICache.scala 55:26]
  reg [52:0] tag1_1; // @[ICache.scala 55:26]
  reg [52:0] tag1_2; // @[ICache.scala 55:26]
  reg [52:0] tag1_3; // @[ICache.scala 55:26]
  reg [52:0] tag1_4; // @[ICache.scala 55:26]
  reg [52:0] tag1_5; // @[ICache.scala 55:26]
  reg [52:0] tag1_6; // @[ICache.scala 55:26]
  reg [52:0] tag1_7; // @[ICache.scala 55:26]
  reg [52:0] tag1_8; // @[ICache.scala 55:26]
  reg [52:0] tag1_9; // @[ICache.scala 55:26]
  reg [52:0] tag1_10; // @[ICache.scala 55:26]
  reg [52:0] tag1_11; // @[ICache.scala 55:26]
  reg [52:0] tag1_12; // @[ICache.scala 55:26]
  reg [52:0] tag1_13; // @[ICache.scala 55:26]
  reg [52:0] tag1_14; // @[ICache.scala 55:26]
  reg [52:0] tag1_15; // @[ICache.scala 55:26]
  reg [52:0] tag1_16; // @[ICache.scala 55:26]
  reg [52:0] tag1_17; // @[ICache.scala 55:26]
  reg [52:0] tag1_18; // @[ICache.scala 55:26]
  reg [52:0] tag1_19; // @[ICache.scala 55:26]
  reg [52:0] tag1_20; // @[ICache.scala 55:26]
  reg [52:0] tag1_21; // @[ICache.scala 55:26]
  reg [52:0] tag1_22; // @[ICache.scala 55:26]
  reg [52:0] tag1_23; // @[ICache.scala 55:26]
  reg [52:0] tag1_24; // @[ICache.scala 55:26]
  reg [52:0] tag1_25; // @[ICache.scala 55:26]
  reg [52:0] tag1_26; // @[ICache.scala 55:26]
  reg [52:0] tag1_27; // @[ICache.scala 55:26]
  reg [52:0] tag1_28; // @[ICache.scala 55:26]
  reg [52:0] tag1_29; // @[ICache.scala 55:26]
  reg [52:0] tag1_30; // @[ICache.scala 55:26]
  reg [52:0] tag1_31; // @[ICache.scala 55:26]
  reg [511:0] block1_0; // @[ICache.scala 56:26]
  reg [511:0] block1_1; // @[ICache.scala 56:26]
  reg [511:0] block1_2; // @[ICache.scala 56:26]
  reg [511:0] block1_3; // @[ICache.scala 56:26]
  reg [511:0] block1_4; // @[ICache.scala 56:26]
  reg [511:0] block1_5; // @[ICache.scala 56:26]
  reg [511:0] block1_6; // @[ICache.scala 56:26]
  reg [511:0] block1_7; // @[ICache.scala 56:26]
  reg [511:0] block1_8; // @[ICache.scala 56:26]
  reg [511:0] block1_9; // @[ICache.scala 56:26]
  reg [511:0] block1_10; // @[ICache.scala 56:26]
  reg [511:0] block1_11; // @[ICache.scala 56:26]
  reg [511:0] block1_12; // @[ICache.scala 56:26]
  reg [511:0] block1_13; // @[ICache.scala 56:26]
  reg [511:0] block1_14; // @[ICache.scala 56:26]
  reg [511:0] block1_15; // @[ICache.scala 56:26]
  reg [511:0] block1_16; // @[ICache.scala 56:26]
  reg [511:0] block1_17; // @[ICache.scala 56:26]
  reg [511:0] block1_18; // @[ICache.scala 56:26]
  reg [511:0] block1_19; // @[ICache.scala 56:26]
  reg [511:0] block1_20; // @[ICache.scala 56:26]
  reg [511:0] block1_21; // @[ICache.scala 56:26]
  reg [511:0] block1_22; // @[ICache.scala 56:26]
  reg [511:0] block1_23; // @[ICache.scala 56:26]
  reg [511:0] block1_24; // @[ICache.scala 56:26]
  reg [511:0] block1_25; // @[ICache.scala 56:26]
  reg [511:0] block1_26; // @[ICache.scala 56:26]
  reg [511:0] block1_27; // @[ICache.scala 56:26]
  reg [511:0] block1_28; // @[ICache.scala 56:26]
  reg [511:0] block1_29; // @[ICache.scala 56:26]
  reg [511:0] block1_30; // @[ICache.scala 56:26]
  reg [511:0] block1_31; // @[ICache.scala 56:26]
  reg  v2_0; // @[ICache.scala 57:26]
  reg  v2_1; // @[ICache.scala 57:26]
  reg  v2_2; // @[ICache.scala 57:26]
  reg  v2_3; // @[ICache.scala 57:26]
  reg  v2_4; // @[ICache.scala 57:26]
  reg  v2_5; // @[ICache.scala 57:26]
  reg  v2_6; // @[ICache.scala 57:26]
  reg  v2_7; // @[ICache.scala 57:26]
  reg  v2_8; // @[ICache.scala 57:26]
  reg  v2_9; // @[ICache.scala 57:26]
  reg  v2_10; // @[ICache.scala 57:26]
  reg  v2_11; // @[ICache.scala 57:26]
  reg  v2_12; // @[ICache.scala 57:26]
  reg  v2_13; // @[ICache.scala 57:26]
  reg  v2_14; // @[ICache.scala 57:26]
  reg  v2_15; // @[ICache.scala 57:26]
  reg  v2_16; // @[ICache.scala 57:26]
  reg  v2_17; // @[ICache.scala 57:26]
  reg  v2_18; // @[ICache.scala 57:26]
  reg  v2_19; // @[ICache.scala 57:26]
  reg  v2_20; // @[ICache.scala 57:26]
  reg  v2_21; // @[ICache.scala 57:26]
  reg  v2_22; // @[ICache.scala 57:26]
  reg  v2_23; // @[ICache.scala 57:26]
  reg  v2_24; // @[ICache.scala 57:26]
  reg  v2_25; // @[ICache.scala 57:26]
  reg  v2_26; // @[ICache.scala 57:26]
  reg  v2_27; // @[ICache.scala 57:26]
  reg  v2_28; // @[ICache.scala 57:26]
  reg  v2_29; // @[ICache.scala 57:26]
  reg  v2_30; // @[ICache.scala 57:26]
  reg  v2_31; // @[ICache.scala 57:26]
  reg  age2_0; // @[ICache.scala 58:26]
  reg  age2_1; // @[ICache.scala 58:26]
  reg  age2_2; // @[ICache.scala 58:26]
  reg  age2_3; // @[ICache.scala 58:26]
  reg  age2_4; // @[ICache.scala 58:26]
  reg  age2_5; // @[ICache.scala 58:26]
  reg  age2_6; // @[ICache.scala 58:26]
  reg  age2_7; // @[ICache.scala 58:26]
  reg  age2_8; // @[ICache.scala 58:26]
  reg  age2_9; // @[ICache.scala 58:26]
  reg  age2_10; // @[ICache.scala 58:26]
  reg  age2_11; // @[ICache.scala 58:26]
  reg  age2_12; // @[ICache.scala 58:26]
  reg  age2_13; // @[ICache.scala 58:26]
  reg  age2_14; // @[ICache.scala 58:26]
  reg  age2_15; // @[ICache.scala 58:26]
  reg  age2_16; // @[ICache.scala 58:26]
  reg  age2_17; // @[ICache.scala 58:26]
  reg  age2_18; // @[ICache.scala 58:26]
  reg  age2_19; // @[ICache.scala 58:26]
  reg  age2_20; // @[ICache.scala 58:26]
  reg  age2_21; // @[ICache.scala 58:26]
  reg  age2_22; // @[ICache.scala 58:26]
  reg  age2_23; // @[ICache.scala 58:26]
  reg  age2_24; // @[ICache.scala 58:26]
  reg  age2_25; // @[ICache.scala 58:26]
  reg  age2_26; // @[ICache.scala 58:26]
  reg  age2_27; // @[ICache.scala 58:26]
  reg  age2_28; // @[ICache.scala 58:26]
  reg  age2_29; // @[ICache.scala 58:26]
  reg  age2_30; // @[ICache.scala 58:26]
  reg  age2_31; // @[ICache.scala 58:26]
  reg [52:0] tag2_0; // @[ICache.scala 59:26]
  reg [52:0] tag2_1; // @[ICache.scala 59:26]
  reg [52:0] tag2_2; // @[ICache.scala 59:26]
  reg [52:0] tag2_3; // @[ICache.scala 59:26]
  reg [52:0] tag2_4; // @[ICache.scala 59:26]
  reg [52:0] tag2_5; // @[ICache.scala 59:26]
  reg [52:0] tag2_6; // @[ICache.scala 59:26]
  reg [52:0] tag2_7; // @[ICache.scala 59:26]
  reg [52:0] tag2_8; // @[ICache.scala 59:26]
  reg [52:0] tag2_9; // @[ICache.scala 59:26]
  reg [52:0] tag2_10; // @[ICache.scala 59:26]
  reg [52:0] tag2_11; // @[ICache.scala 59:26]
  reg [52:0] tag2_12; // @[ICache.scala 59:26]
  reg [52:0] tag2_13; // @[ICache.scala 59:26]
  reg [52:0] tag2_14; // @[ICache.scala 59:26]
  reg [52:0] tag2_15; // @[ICache.scala 59:26]
  reg [52:0] tag2_16; // @[ICache.scala 59:26]
  reg [52:0] tag2_17; // @[ICache.scala 59:26]
  reg [52:0] tag2_18; // @[ICache.scala 59:26]
  reg [52:0] tag2_19; // @[ICache.scala 59:26]
  reg [52:0] tag2_20; // @[ICache.scala 59:26]
  reg [52:0] tag2_21; // @[ICache.scala 59:26]
  reg [52:0] tag2_22; // @[ICache.scala 59:26]
  reg [52:0] tag2_23; // @[ICache.scala 59:26]
  reg [52:0] tag2_24; // @[ICache.scala 59:26]
  reg [52:0] tag2_25; // @[ICache.scala 59:26]
  reg [52:0] tag2_26; // @[ICache.scala 59:26]
  reg [52:0] tag2_27; // @[ICache.scala 59:26]
  reg [52:0] tag2_28; // @[ICache.scala 59:26]
  reg [52:0] tag2_29; // @[ICache.scala 59:26]
  reg [52:0] tag2_30; // @[ICache.scala 59:26]
  reg [52:0] tag2_31; // @[ICache.scala 59:26]
  reg [511:0] block2_0; // @[ICache.scala 60:26]
  reg [511:0] block2_1; // @[ICache.scala 60:26]
  reg [511:0] block2_2; // @[ICache.scala 60:26]
  reg [511:0] block2_3; // @[ICache.scala 60:26]
  reg [511:0] block2_4; // @[ICache.scala 60:26]
  reg [511:0] block2_5; // @[ICache.scala 60:26]
  reg [511:0] block2_6; // @[ICache.scala 60:26]
  reg [511:0] block2_7; // @[ICache.scala 60:26]
  reg [511:0] block2_8; // @[ICache.scala 60:26]
  reg [511:0] block2_9; // @[ICache.scala 60:26]
  reg [511:0] block2_10; // @[ICache.scala 60:26]
  reg [511:0] block2_11; // @[ICache.scala 60:26]
  reg [511:0] block2_12; // @[ICache.scala 60:26]
  reg [511:0] block2_13; // @[ICache.scala 60:26]
  reg [511:0] block2_14; // @[ICache.scala 60:26]
  reg [511:0] block2_15; // @[ICache.scala 60:26]
  reg [511:0] block2_16; // @[ICache.scala 60:26]
  reg [511:0] block2_17; // @[ICache.scala 60:26]
  reg [511:0] block2_18; // @[ICache.scala 60:26]
  reg [511:0] block2_19; // @[ICache.scala 60:26]
  reg [511:0] block2_20; // @[ICache.scala 60:26]
  reg [511:0] block2_21; // @[ICache.scala 60:26]
  reg [511:0] block2_22; // @[ICache.scala 60:26]
  reg [511:0] block2_23; // @[ICache.scala 60:26]
  reg [511:0] block2_24; // @[ICache.scala 60:26]
  reg [511:0] block2_25; // @[ICache.scala 60:26]
  reg [511:0] block2_26; // @[ICache.scala 60:26]
  reg [511:0] block2_27; // @[ICache.scala 60:26]
  reg [511:0] block2_28; // @[ICache.scala 60:26]
  reg [511:0] block2_29; // @[ICache.scala 60:26]
  reg [511:0] block2_30; // @[ICache.scala 60:26]
  reg [511:0] block2_31; // @[ICache.scala 60:26]
  wire [52:0] _GEN_2 = 5'h1 == index_addr ? tag1_1 : tag1_0; // @[ICache.scala 62:28 ICache.scala 62:28]
  wire [52:0] _GEN_3 = 5'h2 == index_addr ? tag1_2 : _GEN_2; // @[ICache.scala 62:28 ICache.scala 62:28]
  wire [52:0] _GEN_4 = 5'h3 == index_addr ? tag1_3 : _GEN_3; // @[ICache.scala 62:28 ICache.scala 62:28]
  wire [52:0] _GEN_5 = 5'h4 == index_addr ? tag1_4 : _GEN_4; // @[ICache.scala 62:28 ICache.scala 62:28]
  wire [52:0] _GEN_6 = 5'h5 == index_addr ? tag1_5 : _GEN_5; // @[ICache.scala 62:28 ICache.scala 62:28]
  wire [52:0] _GEN_7 = 5'h6 == index_addr ? tag1_6 : _GEN_6; // @[ICache.scala 62:28 ICache.scala 62:28]
  wire [52:0] _GEN_8 = 5'h7 == index_addr ? tag1_7 : _GEN_7; // @[ICache.scala 62:28 ICache.scala 62:28]
  wire [52:0] _GEN_9 = 5'h8 == index_addr ? tag1_8 : _GEN_8; // @[ICache.scala 62:28 ICache.scala 62:28]
  wire [52:0] _GEN_10 = 5'h9 == index_addr ? tag1_9 : _GEN_9; // @[ICache.scala 62:28 ICache.scala 62:28]
  wire [52:0] _GEN_11 = 5'ha == index_addr ? tag1_10 : _GEN_10; // @[ICache.scala 62:28 ICache.scala 62:28]
  wire [52:0] _GEN_12 = 5'hb == index_addr ? tag1_11 : _GEN_11; // @[ICache.scala 62:28 ICache.scala 62:28]
  wire [52:0] _GEN_13 = 5'hc == index_addr ? tag1_12 : _GEN_12; // @[ICache.scala 62:28 ICache.scala 62:28]
  wire [52:0] _GEN_14 = 5'hd == index_addr ? tag1_13 : _GEN_13; // @[ICache.scala 62:28 ICache.scala 62:28]
  wire [52:0] _GEN_15 = 5'he == index_addr ? tag1_14 : _GEN_14; // @[ICache.scala 62:28 ICache.scala 62:28]
  wire [52:0] _GEN_16 = 5'hf == index_addr ? tag1_15 : _GEN_15; // @[ICache.scala 62:28 ICache.scala 62:28]
  wire [52:0] _GEN_17 = 5'h10 == index_addr ? tag1_16 : _GEN_16; // @[ICache.scala 62:28 ICache.scala 62:28]
  wire [52:0] _GEN_18 = 5'h11 == index_addr ? tag1_17 : _GEN_17; // @[ICache.scala 62:28 ICache.scala 62:28]
  wire [52:0] _GEN_19 = 5'h12 == index_addr ? tag1_18 : _GEN_18; // @[ICache.scala 62:28 ICache.scala 62:28]
  wire [52:0] _GEN_20 = 5'h13 == index_addr ? tag1_19 : _GEN_19; // @[ICache.scala 62:28 ICache.scala 62:28]
  wire [52:0] _GEN_21 = 5'h14 == index_addr ? tag1_20 : _GEN_20; // @[ICache.scala 62:28 ICache.scala 62:28]
  wire [52:0] _GEN_22 = 5'h15 == index_addr ? tag1_21 : _GEN_21; // @[ICache.scala 62:28 ICache.scala 62:28]
  wire [52:0] _GEN_23 = 5'h16 == index_addr ? tag1_22 : _GEN_22; // @[ICache.scala 62:28 ICache.scala 62:28]
  wire [52:0] _GEN_24 = 5'h17 == index_addr ? tag1_23 : _GEN_23; // @[ICache.scala 62:28 ICache.scala 62:28]
  wire [52:0] _GEN_25 = 5'h18 == index_addr ? tag1_24 : _GEN_24; // @[ICache.scala 62:28 ICache.scala 62:28]
  wire [52:0] _GEN_26 = 5'h19 == index_addr ? tag1_25 : _GEN_25; // @[ICache.scala 62:28 ICache.scala 62:28]
  wire [52:0] _GEN_27 = 5'h1a == index_addr ? tag1_26 : _GEN_26; // @[ICache.scala 62:28 ICache.scala 62:28]
  wire [52:0] _GEN_28 = 5'h1b == index_addr ? tag1_27 : _GEN_27; // @[ICache.scala 62:28 ICache.scala 62:28]
  wire [52:0] _GEN_29 = 5'h1c == index_addr ? tag1_28 : _GEN_28; // @[ICache.scala 62:28 ICache.scala 62:28]
  wire [52:0] _GEN_30 = 5'h1d == index_addr ? tag1_29 : _GEN_29; // @[ICache.scala 62:28 ICache.scala 62:28]
  wire [52:0] _GEN_31 = 5'h1e == index_addr ? tag1_30 : _GEN_30; // @[ICache.scala 62:28 ICache.scala 62:28]
  wire [52:0] _GEN_32 = 5'h1f == index_addr ? tag1_31 : _GEN_31; // @[ICache.scala 62:28 ICache.scala 62:28]
  wire  _GEN_34 = 5'h1 == index_addr ? v1_1 : v1_0; // @[ICache.scala 62:67 ICache.scala 62:67]
  wire  _GEN_35 = 5'h2 == index_addr ? v1_2 : _GEN_34; // @[ICache.scala 62:67 ICache.scala 62:67]
  wire  _GEN_36 = 5'h3 == index_addr ? v1_3 : _GEN_35; // @[ICache.scala 62:67 ICache.scala 62:67]
  wire  _GEN_37 = 5'h4 == index_addr ? v1_4 : _GEN_36; // @[ICache.scala 62:67 ICache.scala 62:67]
  wire  _GEN_38 = 5'h5 == index_addr ? v1_5 : _GEN_37; // @[ICache.scala 62:67 ICache.scala 62:67]
  wire  _GEN_39 = 5'h6 == index_addr ? v1_6 : _GEN_38; // @[ICache.scala 62:67 ICache.scala 62:67]
  wire  _GEN_40 = 5'h7 == index_addr ? v1_7 : _GEN_39; // @[ICache.scala 62:67 ICache.scala 62:67]
  wire  _GEN_41 = 5'h8 == index_addr ? v1_8 : _GEN_40; // @[ICache.scala 62:67 ICache.scala 62:67]
  wire  _GEN_42 = 5'h9 == index_addr ? v1_9 : _GEN_41; // @[ICache.scala 62:67 ICache.scala 62:67]
  wire  _GEN_43 = 5'ha == index_addr ? v1_10 : _GEN_42; // @[ICache.scala 62:67 ICache.scala 62:67]
  wire  _GEN_44 = 5'hb == index_addr ? v1_11 : _GEN_43; // @[ICache.scala 62:67 ICache.scala 62:67]
  wire  _GEN_45 = 5'hc == index_addr ? v1_12 : _GEN_44; // @[ICache.scala 62:67 ICache.scala 62:67]
  wire  _GEN_46 = 5'hd == index_addr ? v1_13 : _GEN_45; // @[ICache.scala 62:67 ICache.scala 62:67]
  wire  _GEN_47 = 5'he == index_addr ? v1_14 : _GEN_46; // @[ICache.scala 62:67 ICache.scala 62:67]
  wire  _GEN_48 = 5'hf == index_addr ? v1_15 : _GEN_47; // @[ICache.scala 62:67 ICache.scala 62:67]
  wire  _GEN_49 = 5'h10 == index_addr ? v1_16 : _GEN_48; // @[ICache.scala 62:67 ICache.scala 62:67]
  wire  _GEN_50 = 5'h11 == index_addr ? v1_17 : _GEN_49; // @[ICache.scala 62:67 ICache.scala 62:67]
  wire  _GEN_51 = 5'h12 == index_addr ? v1_18 : _GEN_50; // @[ICache.scala 62:67 ICache.scala 62:67]
  wire  _GEN_52 = 5'h13 == index_addr ? v1_19 : _GEN_51; // @[ICache.scala 62:67 ICache.scala 62:67]
  wire  _GEN_53 = 5'h14 == index_addr ? v1_20 : _GEN_52; // @[ICache.scala 62:67 ICache.scala 62:67]
  wire  _GEN_54 = 5'h15 == index_addr ? v1_21 : _GEN_53; // @[ICache.scala 62:67 ICache.scala 62:67]
  wire  _GEN_55 = 5'h16 == index_addr ? v1_22 : _GEN_54; // @[ICache.scala 62:67 ICache.scala 62:67]
  wire  _GEN_56 = 5'h17 == index_addr ? v1_23 : _GEN_55; // @[ICache.scala 62:67 ICache.scala 62:67]
  wire  _GEN_57 = 5'h18 == index_addr ? v1_24 : _GEN_56; // @[ICache.scala 62:67 ICache.scala 62:67]
  wire  _GEN_58 = 5'h19 == index_addr ? v1_25 : _GEN_57; // @[ICache.scala 62:67 ICache.scala 62:67]
  wire  _GEN_59 = 5'h1a == index_addr ? v1_26 : _GEN_58; // @[ICache.scala 62:67 ICache.scala 62:67]
  wire  _GEN_60 = 5'h1b == index_addr ? v1_27 : _GEN_59; // @[ICache.scala 62:67 ICache.scala 62:67]
  wire  _GEN_61 = 5'h1c == index_addr ? v1_28 : _GEN_60; // @[ICache.scala 62:67 ICache.scala 62:67]
  wire  _GEN_62 = 5'h1d == index_addr ? v1_29 : _GEN_61; // @[ICache.scala 62:67 ICache.scala 62:67]
  wire  _GEN_63 = 5'h1e == index_addr ? v1_30 : _GEN_62; // @[ICache.scala 62:67 ICache.scala 62:67]
  wire  _GEN_64 = 5'h1f == index_addr ? v1_31 : _GEN_63; // @[ICache.scala 62:67 ICache.scala 62:67]
  wire  hit1 = tag_addr == _GEN_32 & _GEN_64; // @[ICache.scala 62:49]
  wire [52:0] _GEN_66 = 5'h1 == index_addr ? tag2_1 : tag2_0; // @[ICache.scala 63:28 ICache.scala 63:28]
  wire [52:0] _GEN_67 = 5'h2 == index_addr ? tag2_2 : _GEN_66; // @[ICache.scala 63:28 ICache.scala 63:28]
  wire [52:0] _GEN_68 = 5'h3 == index_addr ? tag2_3 : _GEN_67; // @[ICache.scala 63:28 ICache.scala 63:28]
  wire [52:0] _GEN_69 = 5'h4 == index_addr ? tag2_4 : _GEN_68; // @[ICache.scala 63:28 ICache.scala 63:28]
  wire [52:0] _GEN_70 = 5'h5 == index_addr ? tag2_5 : _GEN_69; // @[ICache.scala 63:28 ICache.scala 63:28]
  wire [52:0] _GEN_71 = 5'h6 == index_addr ? tag2_6 : _GEN_70; // @[ICache.scala 63:28 ICache.scala 63:28]
  wire [52:0] _GEN_72 = 5'h7 == index_addr ? tag2_7 : _GEN_71; // @[ICache.scala 63:28 ICache.scala 63:28]
  wire [52:0] _GEN_73 = 5'h8 == index_addr ? tag2_8 : _GEN_72; // @[ICache.scala 63:28 ICache.scala 63:28]
  wire [52:0] _GEN_74 = 5'h9 == index_addr ? tag2_9 : _GEN_73; // @[ICache.scala 63:28 ICache.scala 63:28]
  wire [52:0] _GEN_75 = 5'ha == index_addr ? tag2_10 : _GEN_74; // @[ICache.scala 63:28 ICache.scala 63:28]
  wire [52:0] _GEN_76 = 5'hb == index_addr ? tag2_11 : _GEN_75; // @[ICache.scala 63:28 ICache.scala 63:28]
  wire [52:0] _GEN_77 = 5'hc == index_addr ? tag2_12 : _GEN_76; // @[ICache.scala 63:28 ICache.scala 63:28]
  wire [52:0] _GEN_78 = 5'hd == index_addr ? tag2_13 : _GEN_77; // @[ICache.scala 63:28 ICache.scala 63:28]
  wire [52:0] _GEN_79 = 5'he == index_addr ? tag2_14 : _GEN_78; // @[ICache.scala 63:28 ICache.scala 63:28]
  wire [52:0] _GEN_80 = 5'hf == index_addr ? tag2_15 : _GEN_79; // @[ICache.scala 63:28 ICache.scala 63:28]
  wire [52:0] _GEN_81 = 5'h10 == index_addr ? tag2_16 : _GEN_80; // @[ICache.scala 63:28 ICache.scala 63:28]
  wire [52:0] _GEN_82 = 5'h11 == index_addr ? tag2_17 : _GEN_81; // @[ICache.scala 63:28 ICache.scala 63:28]
  wire [52:0] _GEN_83 = 5'h12 == index_addr ? tag2_18 : _GEN_82; // @[ICache.scala 63:28 ICache.scala 63:28]
  wire [52:0] _GEN_84 = 5'h13 == index_addr ? tag2_19 : _GEN_83; // @[ICache.scala 63:28 ICache.scala 63:28]
  wire [52:0] _GEN_85 = 5'h14 == index_addr ? tag2_20 : _GEN_84; // @[ICache.scala 63:28 ICache.scala 63:28]
  wire [52:0] _GEN_86 = 5'h15 == index_addr ? tag2_21 : _GEN_85; // @[ICache.scala 63:28 ICache.scala 63:28]
  wire [52:0] _GEN_87 = 5'h16 == index_addr ? tag2_22 : _GEN_86; // @[ICache.scala 63:28 ICache.scala 63:28]
  wire [52:0] _GEN_88 = 5'h17 == index_addr ? tag2_23 : _GEN_87; // @[ICache.scala 63:28 ICache.scala 63:28]
  wire [52:0] _GEN_89 = 5'h18 == index_addr ? tag2_24 : _GEN_88; // @[ICache.scala 63:28 ICache.scala 63:28]
  wire [52:0] _GEN_90 = 5'h19 == index_addr ? tag2_25 : _GEN_89; // @[ICache.scala 63:28 ICache.scala 63:28]
  wire [52:0] _GEN_91 = 5'h1a == index_addr ? tag2_26 : _GEN_90; // @[ICache.scala 63:28 ICache.scala 63:28]
  wire [52:0] _GEN_92 = 5'h1b == index_addr ? tag2_27 : _GEN_91; // @[ICache.scala 63:28 ICache.scala 63:28]
  wire [52:0] _GEN_93 = 5'h1c == index_addr ? tag2_28 : _GEN_92; // @[ICache.scala 63:28 ICache.scala 63:28]
  wire [52:0] _GEN_94 = 5'h1d == index_addr ? tag2_29 : _GEN_93; // @[ICache.scala 63:28 ICache.scala 63:28]
  wire [52:0] _GEN_95 = 5'h1e == index_addr ? tag2_30 : _GEN_94; // @[ICache.scala 63:28 ICache.scala 63:28]
  wire [52:0] _GEN_96 = 5'h1f == index_addr ? tag2_31 : _GEN_95; // @[ICache.scala 63:28 ICache.scala 63:28]
  wire  _GEN_98 = 5'h1 == index_addr ? v2_1 : v2_0; // @[ICache.scala 63:67 ICache.scala 63:67]
  wire  _GEN_99 = 5'h2 == index_addr ? v2_2 : _GEN_98; // @[ICache.scala 63:67 ICache.scala 63:67]
  wire  _GEN_100 = 5'h3 == index_addr ? v2_3 : _GEN_99; // @[ICache.scala 63:67 ICache.scala 63:67]
  wire  _GEN_101 = 5'h4 == index_addr ? v2_4 : _GEN_100; // @[ICache.scala 63:67 ICache.scala 63:67]
  wire  _GEN_102 = 5'h5 == index_addr ? v2_5 : _GEN_101; // @[ICache.scala 63:67 ICache.scala 63:67]
  wire  _GEN_103 = 5'h6 == index_addr ? v2_6 : _GEN_102; // @[ICache.scala 63:67 ICache.scala 63:67]
  wire  _GEN_104 = 5'h7 == index_addr ? v2_7 : _GEN_103; // @[ICache.scala 63:67 ICache.scala 63:67]
  wire  _GEN_105 = 5'h8 == index_addr ? v2_8 : _GEN_104; // @[ICache.scala 63:67 ICache.scala 63:67]
  wire  _GEN_106 = 5'h9 == index_addr ? v2_9 : _GEN_105; // @[ICache.scala 63:67 ICache.scala 63:67]
  wire  _GEN_107 = 5'ha == index_addr ? v2_10 : _GEN_106; // @[ICache.scala 63:67 ICache.scala 63:67]
  wire  _GEN_108 = 5'hb == index_addr ? v2_11 : _GEN_107; // @[ICache.scala 63:67 ICache.scala 63:67]
  wire  _GEN_109 = 5'hc == index_addr ? v2_12 : _GEN_108; // @[ICache.scala 63:67 ICache.scala 63:67]
  wire  _GEN_110 = 5'hd == index_addr ? v2_13 : _GEN_109; // @[ICache.scala 63:67 ICache.scala 63:67]
  wire  _GEN_111 = 5'he == index_addr ? v2_14 : _GEN_110; // @[ICache.scala 63:67 ICache.scala 63:67]
  wire  _GEN_112 = 5'hf == index_addr ? v2_15 : _GEN_111; // @[ICache.scala 63:67 ICache.scala 63:67]
  wire  _GEN_113 = 5'h10 == index_addr ? v2_16 : _GEN_112; // @[ICache.scala 63:67 ICache.scala 63:67]
  wire  _GEN_114 = 5'h11 == index_addr ? v2_17 : _GEN_113; // @[ICache.scala 63:67 ICache.scala 63:67]
  wire  _GEN_115 = 5'h12 == index_addr ? v2_18 : _GEN_114; // @[ICache.scala 63:67 ICache.scala 63:67]
  wire  _GEN_116 = 5'h13 == index_addr ? v2_19 : _GEN_115; // @[ICache.scala 63:67 ICache.scala 63:67]
  wire  _GEN_117 = 5'h14 == index_addr ? v2_20 : _GEN_116; // @[ICache.scala 63:67 ICache.scala 63:67]
  wire  _GEN_118 = 5'h15 == index_addr ? v2_21 : _GEN_117; // @[ICache.scala 63:67 ICache.scala 63:67]
  wire  _GEN_119 = 5'h16 == index_addr ? v2_22 : _GEN_118; // @[ICache.scala 63:67 ICache.scala 63:67]
  wire  _GEN_120 = 5'h17 == index_addr ? v2_23 : _GEN_119; // @[ICache.scala 63:67 ICache.scala 63:67]
  wire  _GEN_121 = 5'h18 == index_addr ? v2_24 : _GEN_120; // @[ICache.scala 63:67 ICache.scala 63:67]
  wire  _GEN_122 = 5'h19 == index_addr ? v2_25 : _GEN_121; // @[ICache.scala 63:67 ICache.scala 63:67]
  wire  _GEN_123 = 5'h1a == index_addr ? v2_26 : _GEN_122; // @[ICache.scala 63:67 ICache.scala 63:67]
  wire  _GEN_124 = 5'h1b == index_addr ? v2_27 : _GEN_123; // @[ICache.scala 63:67 ICache.scala 63:67]
  wire  _GEN_125 = 5'h1c == index_addr ? v2_28 : _GEN_124; // @[ICache.scala 63:67 ICache.scala 63:67]
  wire  _GEN_126 = 5'h1d == index_addr ? v2_29 : _GEN_125; // @[ICache.scala 63:67 ICache.scala 63:67]
  wire  _GEN_127 = 5'h1e == index_addr ? v2_30 : _GEN_126; // @[ICache.scala 63:67 ICache.scala 63:67]
  wire  _GEN_128 = 5'h1f == index_addr ? v2_31 : _GEN_127; // @[ICache.scala 63:67 ICache.scala 63:67]
  wire  hit2 = tag_addr == _GEN_96 & _GEN_128; // @[ICache.scala 63:49]
  wire [8:0] _data1_T = {offset_addr, 3'h0}; // @[ICache.scala 64:55]
  wire [511:0] _GEN_130 = 5'h1 == index_addr ? block1_1 : block1_0; // @[ICache.scala 64:39 ICache.scala 64:39]
  wire [511:0] _GEN_131 = 5'h2 == index_addr ? block1_2 : _GEN_130; // @[ICache.scala 64:39 ICache.scala 64:39]
  wire [511:0] _GEN_132 = 5'h3 == index_addr ? block1_3 : _GEN_131; // @[ICache.scala 64:39 ICache.scala 64:39]
  wire [511:0] _GEN_133 = 5'h4 == index_addr ? block1_4 : _GEN_132; // @[ICache.scala 64:39 ICache.scala 64:39]
  wire [511:0] _GEN_134 = 5'h5 == index_addr ? block1_5 : _GEN_133; // @[ICache.scala 64:39 ICache.scala 64:39]
  wire [511:0] _GEN_135 = 5'h6 == index_addr ? block1_6 : _GEN_134; // @[ICache.scala 64:39 ICache.scala 64:39]
  wire [511:0] _GEN_136 = 5'h7 == index_addr ? block1_7 : _GEN_135; // @[ICache.scala 64:39 ICache.scala 64:39]
  wire [511:0] _GEN_137 = 5'h8 == index_addr ? block1_8 : _GEN_136; // @[ICache.scala 64:39 ICache.scala 64:39]
  wire [511:0] _GEN_138 = 5'h9 == index_addr ? block1_9 : _GEN_137; // @[ICache.scala 64:39 ICache.scala 64:39]
  wire [511:0] _GEN_139 = 5'ha == index_addr ? block1_10 : _GEN_138; // @[ICache.scala 64:39 ICache.scala 64:39]
  wire [511:0] _GEN_140 = 5'hb == index_addr ? block1_11 : _GEN_139; // @[ICache.scala 64:39 ICache.scala 64:39]
  wire [511:0] _GEN_141 = 5'hc == index_addr ? block1_12 : _GEN_140; // @[ICache.scala 64:39 ICache.scala 64:39]
  wire [511:0] _GEN_142 = 5'hd == index_addr ? block1_13 : _GEN_141; // @[ICache.scala 64:39 ICache.scala 64:39]
  wire [511:0] _GEN_143 = 5'he == index_addr ? block1_14 : _GEN_142; // @[ICache.scala 64:39 ICache.scala 64:39]
  wire [511:0] _GEN_144 = 5'hf == index_addr ? block1_15 : _GEN_143; // @[ICache.scala 64:39 ICache.scala 64:39]
  wire [511:0] _GEN_145 = 5'h10 == index_addr ? block1_16 : _GEN_144; // @[ICache.scala 64:39 ICache.scala 64:39]
  wire [511:0] _GEN_146 = 5'h11 == index_addr ? block1_17 : _GEN_145; // @[ICache.scala 64:39 ICache.scala 64:39]
  wire [511:0] _GEN_147 = 5'h12 == index_addr ? block1_18 : _GEN_146; // @[ICache.scala 64:39 ICache.scala 64:39]
  wire [511:0] _GEN_148 = 5'h13 == index_addr ? block1_19 : _GEN_147; // @[ICache.scala 64:39 ICache.scala 64:39]
  wire [511:0] _GEN_149 = 5'h14 == index_addr ? block1_20 : _GEN_148; // @[ICache.scala 64:39 ICache.scala 64:39]
  wire [511:0] _GEN_150 = 5'h15 == index_addr ? block1_21 : _GEN_149; // @[ICache.scala 64:39 ICache.scala 64:39]
  wire [511:0] _GEN_151 = 5'h16 == index_addr ? block1_22 : _GEN_150; // @[ICache.scala 64:39 ICache.scala 64:39]
  wire [511:0] _GEN_152 = 5'h17 == index_addr ? block1_23 : _GEN_151; // @[ICache.scala 64:39 ICache.scala 64:39]
  wire [511:0] _GEN_153 = 5'h18 == index_addr ? block1_24 : _GEN_152; // @[ICache.scala 64:39 ICache.scala 64:39]
  wire [511:0] _GEN_154 = 5'h19 == index_addr ? block1_25 : _GEN_153; // @[ICache.scala 64:39 ICache.scala 64:39]
  wire [511:0] _GEN_155 = 5'h1a == index_addr ? block1_26 : _GEN_154; // @[ICache.scala 64:39 ICache.scala 64:39]
  wire [511:0] _GEN_156 = 5'h1b == index_addr ? block1_27 : _GEN_155; // @[ICache.scala 64:39 ICache.scala 64:39]
  wire [511:0] _GEN_157 = 5'h1c == index_addr ? block1_28 : _GEN_156; // @[ICache.scala 64:39 ICache.scala 64:39]
  wire [511:0] _GEN_158 = 5'h1d == index_addr ? block1_29 : _GEN_157; // @[ICache.scala 64:39 ICache.scala 64:39]
  wire [511:0] _GEN_159 = 5'h1e == index_addr ? block1_30 : _GEN_158; // @[ICache.scala 64:39 ICache.scala 64:39]
  wire [511:0] _GEN_160 = 5'h1f == index_addr ? block1_31 : _GEN_159; // @[ICache.scala 64:39 ICache.scala 64:39]
  wire [511:0] _data1_T_1 = _GEN_160 >> _data1_T; // @[ICache.scala 64:39]
  wire [31:0] data1 = _data1_T_1[31:0]; // @[ICache.scala 64:61]
  wire [511:0] _GEN_162 = 5'h1 == index_addr ? block2_1 : block2_0; // @[ICache.scala 65:39 ICache.scala 65:39]
  wire [511:0] _GEN_163 = 5'h2 == index_addr ? block2_2 : _GEN_162; // @[ICache.scala 65:39 ICache.scala 65:39]
  wire [511:0] _GEN_164 = 5'h3 == index_addr ? block2_3 : _GEN_163; // @[ICache.scala 65:39 ICache.scala 65:39]
  wire [511:0] _GEN_165 = 5'h4 == index_addr ? block2_4 : _GEN_164; // @[ICache.scala 65:39 ICache.scala 65:39]
  wire [511:0] _GEN_166 = 5'h5 == index_addr ? block2_5 : _GEN_165; // @[ICache.scala 65:39 ICache.scala 65:39]
  wire [511:0] _GEN_167 = 5'h6 == index_addr ? block2_6 : _GEN_166; // @[ICache.scala 65:39 ICache.scala 65:39]
  wire [511:0] _GEN_168 = 5'h7 == index_addr ? block2_7 : _GEN_167; // @[ICache.scala 65:39 ICache.scala 65:39]
  wire [511:0] _GEN_169 = 5'h8 == index_addr ? block2_8 : _GEN_168; // @[ICache.scala 65:39 ICache.scala 65:39]
  wire [511:0] _GEN_170 = 5'h9 == index_addr ? block2_9 : _GEN_169; // @[ICache.scala 65:39 ICache.scala 65:39]
  wire [511:0] _GEN_171 = 5'ha == index_addr ? block2_10 : _GEN_170; // @[ICache.scala 65:39 ICache.scala 65:39]
  wire [511:0] _GEN_172 = 5'hb == index_addr ? block2_11 : _GEN_171; // @[ICache.scala 65:39 ICache.scala 65:39]
  wire [511:0] _GEN_173 = 5'hc == index_addr ? block2_12 : _GEN_172; // @[ICache.scala 65:39 ICache.scala 65:39]
  wire [511:0] _GEN_174 = 5'hd == index_addr ? block2_13 : _GEN_173; // @[ICache.scala 65:39 ICache.scala 65:39]
  wire [511:0] _GEN_175 = 5'he == index_addr ? block2_14 : _GEN_174; // @[ICache.scala 65:39 ICache.scala 65:39]
  wire [511:0] _GEN_176 = 5'hf == index_addr ? block2_15 : _GEN_175; // @[ICache.scala 65:39 ICache.scala 65:39]
  wire [511:0] _GEN_177 = 5'h10 == index_addr ? block2_16 : _GEN_176; // @[ICache.scala 65:39 ICache.scala 65:39]
  wire [511:0] _GEN_178 = 5'h11 == index_addr ? block2_17 : _GEN_177; // @[ICache.scala 65:39 ICache.scala 65:39]
  wire [511:0] _GEN_179 = 5'h12 == index_addr ? block2_18 : _GEN_178; // @[ICache.scala 65:39 ICache.scala 65:39]
  wire [511:0] _GEN_180 = 5'h13 == index_addr ? block2_19 : _GEN_179; // @[ICache.scala 65:39 ICache.scala 65:39]
  wire [511:0] _GEN_181 = 5'h14 == index_addr ? block2_20 : _GEN_180; // @[ICache.scala 65:39 ICache.scala 65:39]
  wire [511:0] _GEN_182 = 5'h15 == index_addr ? block2_21 : _GEN_181; // @[ICache.scala 65:39 ICache.scala 65:39]
  wire [511:0] _GEN_183 = 5'h16 == index_addr ? block2_22 : _GEN_182; // @[ICache.scala 65:39 ICache.scala 65:39]
  wire [511:0] _GEN_184 = 5'h17 == index_addr ? block2_23 : _GEN_183; // @[ICache.scala 65:39 ICache.scala 65:39]
  wire [511:0] _GEN_185 = 5'h18 == index_addr ? block2_24 : _GEN_184; // @[ICache.scala 65:39 ICache.scala 65:39]
  wire [511:0] _GEN_186 = 5'h19 == index_addr ? block2_25 : _GEN_185; // @[ICache.scala 65:39 ICache.scala 65:39]
  wire [511:0] _GEN_187 = 5'h1a == index_addr ? block2_26 : _GEN_186; // @[ICache.scala 65:39 ICache.scala 65:39]
  wire [511:0] _GEN_188 = 5'h1b == index_addr ? block2_27 : _GEN_187; // @[ICache.scala 65:39 ICache.scala 65:39]
  wire [511:0] _GEN_189 = 5'h1c == index_addr ? block2_28 : _GEN_188; // @[ICache.scala 65:39 ICache.scala 65:39]
  wire [511:0] _GEN_190 = 5'h1d == index_addr ? block2_29 : _GEN_189; // @[ICache.scala 65:39 ICache.scala 65:39]
  wire [511:0] _GEN_191 = 5'h1e == index_addr ? block2_30 : _GEN_190; // @[ICache.scala 65:39 ICache.scala 65:39]
  wire [511:0] _GEN_192 = 5'h1f == index_addr ? block2_31 : _GEN_191; // @[ICache.scala 65:39 ICache.scala 65:39]
  wire [511:0] _data2_T_1 = _GEN_192 >> _data1_T; // @[ICache.scala 65:39]
  wire [31:0] data2 = _data2_T_1[31:0]; // @[ICache.scala 65:61]
  wire  hit = hit1 | hit2; // @[ICache.scala 67:24]
  wire [31:0] _data_T = hit1 ? data1 : 32'h0; // @[ICache.scala 68:39]
  wire  _age1_T = hit1 ^ hit2; // @[ICache.scala 71:34]
  wire  _GEN_194 = 5'h1 == index_addr ? age1_1 : age1_0; // @[ICache.scala 71:28 ICache.scala 71:28]
  wire  _GEN_195 = 5'h2 == index_addr ? age1_2 : _GEN_194; // @[ICache.scala 71:28 ICache.scala 71:28]
  wire  _GEN_196 = 5'h3 == index_addr ? age1_3 : _GEN_195; // @[ICache.scala 71:28 ICache.scala 71:28]
  wire  _GEN_197 = 5'h4 == index_addr ? age1_4 : _GEN_196; // @[ICache.scala 71:28 ICache.scala 71:28]
  wire  _GEN_198 = 5'h5 == index_addr ? age1_5 : _GEN_197; // @[ICache.scala 71:28 ICache.scala 71:28]
  wire  _GEN_199 = 5'h6 == index_addr ? age1_6 : _GEN_198; // @[ICache.scala 71:28 ICache.scala 71:28]
  wire  _GEN_200 = 5'h7 == index_addr ? age1_7 : _GEN_199; // @[ICache.scala 71:28 ICache.scala 71:28]
  wire  _GEN_201 = 5'h8 == index_addr ? age1_8 : _GEN_200; // @[ICache.scala 71:28 ICache.scala 71:28]
  wire  _GEN_202 = 5'h9 == index_addr ? age1_9 : _GEN_201; // @[ICache.scala 71:28 ICache.scala 71:28]
  wire  _GEN_203 = 5'ha == index_addr ? age1_10 : _GEN_202; // @[ICache.scala 71:28 ICache.scala 71:28]
  wire  _GEN_204 = 5'hb == index_addr ? age1_11 : _GEN_203; // @[ICache.scala 71:28 ICache.scala 71:28]
  wire  _GEN_205 = 5'hc == index_addr ? age1_12 : _GEN_204; // @[ICache.scala 71:28 ICache.scala 71:28]
  wire  _GEN_206 = 5'hd == index_addr ? age1_13 : _GEN_205; // @[ICache.scala 71:28 ICache.scala 71:28]
  wire  _GEN_207 = 5'he == index_addr ? age1_14 : _GEN_206; // @[ICache.scala 71:28 ICache.scala 71:28]
  wire  _GEN_208 = 5'hf == index_addr ? age1_15 : _GEN_207; // @[ICache.scala 71:28 ICache.scala 71:28]
  wire  _GEN_209 = 5'h10 == index_addr ? age1_16 : _GEN_208; // @[ICache.scala 71:28 ICache.scala 71:28]
  wire  _GEN_210 = 5'h11 == index_addr ? age1_17 : _GEN_209; // @[ICache.scala 71:28 ICache.scala 71:28]
  wire  _GEN_211 = 5'h12 == index_addr ? age1_18 : _GEN_210; // @[ICache.scala 71:28 ICache.scala 71:28]
  wire  _GEN_212 = 5'h13 == index_addr ? age1_19 : _GEN_211; // @[ICache.scala 71:28 ICache.scala 71:28]
  wire  _GEN_213 = 5'h14 == index_addr ? age1_20 : _GEN_212; // @[ICache.scala 71:28 ICache.scala 71:28]
  wire  _GEN_214 = 5'h15 == index_addr ? age1_21 : _GEN_213; // @[ICache.scala 71:28 ICache.scala 71:28]
  wire  _GEN_215 = 5'h16 == index_addr ? age1_22 : _GEN_214; // @[ICache.scala 71:28 ICache.scala 71:28]
  wire  _GEN_216 = 5'h17 == index_addr ? age1_23 : _GEN_215; // @[ICache.scala 71:28 ICache.scala 71:28]
  wire  _GEN_217 = 5'h18 == index_addr ? age1_24 : _GEN_216; // @[ICache.scala 71:28 ICache.scala 71:28]
  wire  _GEN_218 = 5'h19 == index_addr ? age1_25 : _GEN_217; // @[ICache.scala 71:28 ICache.scala 71:28]
  wire  _GEN_219 = 5'h1a == index_addr ? age1_26 : _GEN_218; // @[ICache.scala 71:28 ICache.scala 71:28]
  wire  _GEN_220 = 5'h1b == index_addr ? age1_27 : _GEN_219; // @[ICache.scala 71:28 ICache.scala 71:28]
  wire  _GEN_221 = 5'h1c == index_addr ? age1_28 : _GEN_220; // @[ICache.scala 71:28 ICache.scala 71:28]
  wire  _GEN_222 = 5'h1d == index_addr ? age1_29 : _GEN_221; // @[ICache.scala 71:28 ICache.scala 71:28]
  wire  _GEN_223 = 5'h1e == index_addr ? age1_30 : _GEN_222; // @[ICache.scala 71:28 ICache.scala 71:28]
  wire  _GEN_224 = 5'h1f == index_addr ? age1_31 : _GEN_223; // @[ICache.scala 71:28 ICache.scala 71:28]
  wire  _GEN_258 = 5'h1 == index_addr ? age2_1 : age2_0; // @[ICache.scala 72:28 ICache.scala 72:28]
  wire  _GEN_259 = 5'h2 == index_addr ? age2_2 : _GEN_258; // @[ICache.scala 72:28 ICache.scala 72:28]
  wire  _GEN_260 = 5'h3 == index_addr ? age2_3 : _GEN_259; // @[ICache.scala 72:28 ICache.scala 72:28]
  wire  _GEN_261 = 5'h4 == index_addr ? age2_4 : _GEN_260; // @[ICache.scala 72:28 ICache.scala 72:28]
  wire  _GEN_262 = 5'h5 == index_addr ? age2_5 : _GEN_261; // @[ICache.scala 72:28 ICache.scala 72:28]
  wire  _GEN_263 = 5'h6 == index_addr ? age2_6 : _GEN_262; // @[ICache.scala 72:28 ICache.scala 72:28]
  wire  _GEN_264 = 5'h7 == index_addr ? age2_7 : _GEN_263; // @[ICache.scala 72:28 ICache.scala 72:28]
  wire  _GEN_265 = 5'h8 == index_addr ? age2_8 : _GEN_264; // @[ICache.scala 72:28 ICache.scala 72:28]
  wire  _GEN_266 = 5'h9 == index_addr ? age2_9 : _GEN_265; // @[ICache.scala 72:28 ICache.scala 72:28]
  wire  _GEN_267 = 5'ha == index_addr ? age2_10 : _GEN_266; // @[ICache.scala 72:28 ICache.scala 72:28]
  wire  _GEN_268 = 5'hb == index_addr ? age2_11 : _GEN_267; // @[ICache.scala 72:28 ICache.scala 72:28]
  wire  _GEN_269 = 5'hc == index_addr ? age2_12 : _GEN_268; // @[ICache.scala 72:28 ICache.scala 72:28]
  wire  _GEN_270 = 5'hd == index_addr ? age2_13 : _GEN_269; // @[ICache.scala 72:28 ICache.scala 72:28]
  wire  _GEN_271 = 5'he == index_addr ? age2_14 : _GEN_270; // @[ICache.scala 72:28 ICache.scala 72:28]
  wire  _GEN_272 = 5'hf == index_addr ? age2_15 : _GEN_271; // @[ICache.scala 72:28 ICache.scala 72:28]
  wire  _GEN_273 = 5'h10 == index_addr ? age2_16 : _GEN_272; // @[ICache.scala 72:28 ICache.scala 72:28]
  wire  _GEN_274 = 5'h11 == index_addr ? age2_17 : _GEN_273; // @[ICache.scala 72:28 ICache.scala 72:28]
  wire  _GEN_275 = 5'h12 == index_addr ? age2_18 : _GEN_274; // @[ICache.scala 72:28 ICache.scala 72:28]
  wire  _GEN_276 = 5'h13 == index_addr ? age2_19 : _GEN_275; // @[ICache.scala 72:28 ICache.scala 72:28]
  wire  _GEN_277 = 5'h14 == index_addr ? age2_20 : _GEN_276; // @[ICache.scala 72:28 ICache.scala 72:28]
  wire  _GEN_278 = 5'h15 == index_addr ? age2_21 : _GEN_277; // @[ICache.scala 72:28 ICache.scala 72:28]
  wire  _GEN_279 = 5'h16 == index_addr ? age2_22 : _GEN_278; // @[ICache.scala 72:28 ICache.scala 72:28]
  wire  _GEN_280 = 5'h17 == index_addr ? age2_23 : _GEN_279; // @[ICache.scala 72:28 ICache.scala 72:28]
  wire  _GEN_281 = 5'h18 == index_addr ? age2_24 : _GEN_280; // @[ICache.scala 72:28 ICache.scala 72:28]
  wire  _GEN_282 = 5'h19 == index_addr ? age2_25 : _GEN_281; // @[ICache.scala 72:28 ICache.scala 72:28]
  wire  _GEN_283 = 5'h1a == index_addr ? age2_26 : _GEN_282; // @[ICache.scala 72:28 ICache.scala 72:28]
  wire  _GEN_284 = 5'h1b == index_addr ? age2_27 : _GEN_283; // @[ICache.scala 72:28 ICache.scala 72:28]
  wire  _GEN_285 = 5'h1c == index_addr ? age2_28 : _GEN_284; // @[ICache.scala 72:28 ICache.scala 72:28]
  wire  _GEN_286 = 5'h1d == index_addr ? age2_29 : _GEN_285; // @[ICache.scala 72:28 ICache.scala 72:28]
  wire  _GEN_287 = 5'h1e == index_addr ? age2_30 : _GEN_286; // @[ICache.scala 72:28 ICache.scala 72:28]
  wire  _GEN_288 = 5'h1f == index_addr ? age2_31 : _GEN_287; // @[ICache.scala 72:28 ICache.scala 72:28]
  reg [1:0] state; // @[ICache.scala 75:24]
  reg  not_en_yet; // @[ICache.scala 78:30]
  wire  _not_en_yet_T = io_imem_en ? 1'h0 : not_en_yet; // @[ICache.scala 79:27]
  reg [4:0] fence_cnt; // @[ICache.scala 84:28]
  wire  _T = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_4 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_5 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_6 = fence_cnt == 5'h1f; // @[ICache.scala 94:28]
  wire [1:0] _GEN_324 = fence_cnt == 5'h1f ? 2'h3 : state; // @[ICache.scala 94:53 ICache.scala 94:60 ICache.scala 75:24]
  wire  _T_7 = 2'h3 == state; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_325 = _T_6 ? 2'h0 : state; // @[ICache.scala 97:53 ICache.scala 97:60 ICache.scala 75:24]
  wire [1:0] _GEN_326 = _T_7 ? _GEN_325 : state; // @[Conditional.scala 39:67 ICache.scala 75:24]
  wire  _io_axi_req_T = state == 2'h1; // @[ICache.scala 102:28]
  wire [1:0] age = {_GEN_288,_GEN_224}; // @[Cat.scala 30:58]
  wire  updateway2 = age == 2'h1; // @[ICache.scala 107:26]
  wire  updateway1 = ~updateway2; // @[ICache.scala 108:22]
  wire  update = _io_axi_req_T & io_axi_valid; // @[ICache.scala 109:33]
  wire  _block1_T = update & updateway1; // @[ICache.scala 110:40]
  wire  _GEN_394 = 5'h0 == index_addr ? _block1_T | _GEN_64 : v1_0; // @[ICache.scala 112:26 ICache.scala 112:26 ICache.scala 53:26]
  wire  _GEN_395 = 5'h1 == index_addr ? _block1_T | _GEN_64 : v1_1; // @[ICache.scala 112:26 ICache.scala 112:26 ICache.scala 53:26]
  wire  _GEN_396 = 5'h2 == index_addr ? _block1_T | _GEN_64 : v1_2; // @[ICache.scala 112:26 ICache.scala 112:26 ICache.scala 53:26]
  wire  _GEN_397 = 5'h3 == index_addr ? _block1_T | _GEN_64 : v1_3; // @[ICache.scala 112:26 ICache.scala 112:26 ICache.scala 53:26]
  wire  _GEN_398 = 5'h4 == index_addr ? _block1_T | _GEN_64 : v1_4; // @[ICache.scala 112:26 ICache.scala 112:26 ICache.scala 53:26]
  wire  _GEN_399 = 5'h5 == index_addr ? _block1_T | _GEN_64 : v1_5; // @[ICache.scala 112:26 ICache.scala 112:26 ICache.scala 53:26]
  wire  _GEN_400 = 5'h6 == index_addr ? _block1_T | _GEN_64 : v1_6; // @[ICache.scala 112:26 ICache.scala 112:26 ICache.scala 53:26]
  wire  _GEN_401 = 5'h7 == index_addr ? _block1_T | _GEN_64 : v1_7; // @[ICache.scala 112:26 ICache.scala 112:26 ICache.scala 53:26]
  wire  _GEN_402 = 5'h8 == index_addr ? _block1_T | _GEN_64 : v1_8; // @[ICache.scala 112:26 ICache.scala 112:26 ICache.scala 53:26]
  wire  _GEN_403 = 5'h9 == index_addr ? _block1_T | _GEN_64 : v1_9; // @[ICache.scala 112:26 ICache.scala 112:26 ICache.scala 53:26]
  wire  _GEN_404 = 5'ha == index_addr ? _block1_T | _GEN_64 : v1_10; // @[ICache.scala 112:26 ICache.scala 112:26 ICache.scala 53:26]
  wire  _GEN_405 = 5'hb == index_addr ? _block1_T | _GEN_64 : v1_11; // @[ICache.scala 112:26 ICache.scala 112:26 ICache.scala 53:26]
  wire  _GEN_406 = 5'hc == index_addr ? _block1_T | _GEN_64 : v1_12; // @[ICache.scala 112:26 ICache.scala 112:26 ICache.scala 53:26]
  wire  _GEN_407 = 5'hd == index_addr ? _block1_T | _GEN_64 : v1_13; // @[ICache.scala 112:26 ICache.scala 112:26 ICache.scala 53:26]
  wire  _GEN_408 = 5'he == index_addr ? _block1_T | _GEN_64 : v1_14; // @[ICache.scala 112:26 ICache.scala 112:26 ICache.scala 53:26]
  wire  _GEN_409 = 5'hf == index_addr ? _block1_T | _GEN_64 : v1_15; // @[ICache.scala 112:26 ICache.scala 112:26 ICache.scala 53:26]
  wire  _GEN_410 = 5'h10 == index_addr ? _block1_T | _GEN_64 : v1_16; // @[ICache.scala 112:26 ICache.scala 112:26 ICache.scala 53:26]
  wire  _GEN_411 = 5'h11 == index_addr ? _block1_T | _GEN_64 : v1_17; // @[ICache.scala 112:26 ICache.scala 112:26 ICache.scala 53:26]
  wire  _GEN_412 = 5'h12 == index_addr ? _block1_T | _GEN_64 : v1_18; // @[ICache.scala 112:26 ICache.scala 112:26 ICache.scala 53:26]
  wire  _GEN_413 = 5'h13 == index_addr ? _block1_T | _GEN_64 : v1_19; // @[ICache.scala 112:26 ICache.scala 112:26 ICache.scala 53:26]
  wire  _GEN_414 = 5'h14 == index_addr ? _block1_T | _GEN_64 : v1_20; // @[ICache.scala 112:26 ICache.scala 112:26 ICache.scala 53:26]
  wire  _GEN_415 = 5'h15 == index_addr ? _block1_T | _GEN_64 : v1_21; // @[ICache.scala 112:26 ICache.scala 112:26 ICache.scala 53:26]
  wire  _GEN_416 = 5'h16 == index_addr ? _block1_T | _GEN_64 : v1_22; // @[ICache.scala 112:26 ICache.scala 112:26 ICache.scala 53:26]
  wire  _GEN_417 = 5'h17 == index_addr ? _block1_T | _GEN_64 : v1_23; // @[ICache.scala 112:26 ICache.scala 112:26 ICache.scala 53:26]
  wire  _GEN_418 = 5'h18 == index_addr ? _block1_T | _GEN_64 : v1_24; // @[ICache.scala 112:26 ICache.scala 112:26 ICache.scala 53:26]
  wire  _GEN_419 = 5'h19 == index_addr ? _block1_T | _GEN_64 : v1_25; // @[ICache.scala 112:26 ICache.scala 112:26 ICache.scala 53:26]
  wire  _GEN_420 = 5'h1a == index_addr ? _block1_T | _GEN_64 : v1_26; // @[ICache.scala 112:26 ICache.scala 112:26 ICache.scala 53:26]
  wire  _GEN_421 = 5'h1b == index_addr ? _block1_T | _GEN_64 : v1_27; // @[ICache.scala 112:26 ICache.scala 112:26 ICache.scala 53:26]
  wire  _GEN_422 = 5'h1c == index_addr ? _block1_T | _GEN_64 : v1_28; // @[ICache.scala 112:26 ICache.scala 112:26 ICache.scala 53:26]
  wire  _GEN_423 = 5'h1d == index_addr ? _block1_T | _GEN_64 : v1_29; // @[ICache.scala 112:26 ICache.scala 112:26 ICache.scala 53:26]
  wire  _GEN_424 = 5'h1e == index_addr ? _block1_T | _GEN_64 : v1_30; // @[ICache.scala 112:26 ICache.scala 112:26 ICache.scala 53:26]
  wire  _GEN_425 = 5'h1f == index_addr ? _block1_T | _GEN_64 : v1_31; // @[ICache.scala 112:26 ICache.scala 112:26 ICache.scala 53:26]
  wire  _block2_T = update & updateway2; // @[ICache.scala 113:40]
  wire  _GEN_490 = 5'h0 == index_addr ? _block2_T | _GEN_128 : v2_0; // @[ICache.scala 115:26 ICache.scala 115:26 ICache.scala 57:26]
  wire  _GEN_491 = 5'h1 == index_addr ? _block2_T | _GEN_128 : v2_1; // @[ICache.scala 115:26 ICache.scala 115:26 ICache.scala 57:26]
  wire  _GEN_492 = 5'h2 == index_addr ? _block2_T | _GEN_128 : v2_2; // @[ICache.scala 115:26 ICache.scala 115:26 ICache.scala 57:26]
  wire  _GEN_493 = 5'h3 == index_addr ? _block2_T | _GEN_128 : v2_3; // @[ICache.scala 115:26 ICache.scala 115:26 ICache.scala 57:26]
  wire  _GEN_494 = 5'h4 == index_addr ? _block2_T | _GEN_128 : v2_4; // @[ICache.scala 115:26 ICache.scala 115:26 ICache.scala 57:26]
  wire  _GEN_495 = 5'h5 == index_addr ? _block2_T | _GEN_128 : v2_5; // @[ICache.scala 115:26 ICache.scala 115:26 ICache.scala 57:26]
  wire  _GEN_496 = 5'h6 == index_addr ? _block2_T | _GEN_128 : v2_6; // @[ICache.scala 115:26 ICache.scala 115:26 ICache.scala 57:26]
  wire  _GEN_497 = 5'h7 == index_addr ? _block2_T | _GEN_128 : v2_7; // @[ICache.scala 115:26 ICache.scala 115:26 ICache.scala 57:26]
  wire  _GEN_498 = 5'h8 == index_addr ? _block2_T | _GEN_128 : v2_8; // @[ICache.scala 115:26 ICache.scala 115:26 ICache.scala 57:26]
  wire  _GEN_499 = 5'h9 == index_addr ? _block2_T | _GEN_128 : v2_9; // @[ICache.scala 115:26 ICache.scala 115:26 ICache.scala 57:26]
  wire  _GEN_500 = 5'ha == index_addr ? _block2_T | _GEN_128 : v2_10; // @[ICache.scala 115:26 ICache.scala 115:26 ICache.scala 57:26]
  wire  _GEN_501 = 5'hb == index_addr ? _block2_T | _GEN_128 : v2_11; // @[ICache.scala 115:26 ICache.scala 115:26 ICache.scala 57:26]
  wire  _GEN_502 = 5'hc == index_addr ? _block2_T | _GEN_128 : v2_12; // @[ICache.scala 115:26 ICache.scala 115:26 ICache.scala 57:26]
  wire  _GEN_503 = 5'hd == index_addr ? _block2_T | _GEN_128 : v2_13; // @[ICache.scala 115:26 ICache.scala 115:26 ICache.scala 57:26]
  wire  _GEN_504 = 5'he == index_addr ? _block2_T | _GEN_128 : v2_14; // @[ICache.scala 115:26 ICache.scala 115:26 ICache.scala 57:26]
  wire  _GEN_505 = 5'hf == index_addr ? _block2_T | _GEN_128 : v2_15; // @[ICache.scala 115:26 ICache.scala 115:26 ICache.scala 57:26]
  wire  _GEN_506 = 5'h10 == index_addr ? _block2_T | _GEN_128 : v2_16; // @[ICache.scala 115:26 ICache.scala 115:26 ICache.scala 57:26]
  wire  _GEN_507 = 5'h11 == index_addr ? _block2_T | _GEN_128 : v2_17; // @[ICache.scala 115:26 ICache.scala 115:26 ICache.scala 57:26]
  wire  _GEN_508 = 5'h12 == index_addr ? _block2_T | _GEN_128 : v2_18; // @[ICache.scala 115:26 ICache.scala 115:26 ICache.scala 57:26]
  wire  _GEN_509 = 5'h13 == index_addr ? _block2_T | _GEN_128 : v2_19; // @[ICache.scala 115:26 ICache.scala 115:26 ICache.scala 57:26]
  wire  _GEN_510 = 5'h14 == index_addr ? _block2_T | _GEN_128 : v2_20; // @[ICache.scala 115:26 ICache.scala 115:26 ICache.scala 57:26]
  wire  _GEN_511 = 5'h15 == index_addr ? _block2_T | _GEN_128 : v2_21; // @[ICache.scala 115:26 ICache.scala 115:26 ICache.scala 57:26]
  wire  _GEN_512 = 5'h16 == index_addr ? _block2_T | _GEN_128 : v2_22; // @[ICache.scala 115:26 ICache.scala 115:26 ICache.scala 57:26]
  wire  _GEN_513 = 5'h17 == index_addr ? _block2_T | _GEN_128 : v2_23; // @[ICache.scala 115:26 ICache.scala 115:26 ICache.scala 57:26]
  wire  _GEN_514 = 5'h18 == index_addr ? _block2_T | _GEN_128 : v2_24; // @[ICache.scala 115:26 ICache.scala 115:26 ICache.scala 57:26]
  wire  _GEN_515 = 5'h19 == index_addr ? _block2_T | _GEN_128 : v2_25; // @[ICache.scala 115:26 ICache.scala 115:26 ICache.scala 57:26]
  wire  _GEN_516 = 5'h1a == index_addr ? _block2_T | _GEN_128 : v2_26; // @[ICache.scala 115:26 ICache.scala 115:26 ICache.scala 57:26]
  wire  _GEN_517 = 5'h1b == index_addr ? _block2_T | _GEN_128 : v2_27; // @[ICache.scala 115:26 ICache.scala 115:26 ICache.scala 57:26]
  wire  _GEN_518 = 5'h1c == index_addr ? _block2_T | _GEN_128 : v2_28; // @[ICache.scala 115:26 ICache.scala 115:26 ICache.scala 57:26]
  wire  _GEN_519 = 5'h1d == index_addr ? _block2_T | _GEN_128 : v2_29; // @[ICache.scala 115:26 ICache.scala 115:26 ICache.scala 57:26]
  wire  _GEN_520 = 5'h1e == index_addr ? _block2_T | _GEN_128 : v2_30; // @[ICache.scala 115:26 ICache.scala 115:26 ICache.scala 57:26]
  wire  _GEN_521 = 5'h1f == index_addr ? _block2_T | _GEN_128 : v2_31; // @[ICache.scala 115:26 ICache.scala 115:26 ICache.scala 57:26]
  wire  _T_9 = state == 2'h2; // @[ICache.scala 117:16]
  wire  _GEN_779 = 5'h0 == index_addr; // @[ICache.scala 118:53 ICache.scala 118:53]
  wire  _GEN_780 = 5'h1 == index_addr; // @[ICache.scala 118:53 ICache.scala 118:53]
  wire  _GEN_781 = 5'h2 == index_addr; // @[ICache.scala 118:53 ICache.scala 118:53]
  wire  _GEN_782 = 5'h3 == index_addr; // @[ICache.scala 118:53 ICache.scala 118:53]
  wire  _GEN_783 = 5'h4 == index_addr; // @[ICache.scala 118:53 ICache.scala 118:53]
  wire  _GEN_784 = 5'h5 == index_addr; // @[ICache.scala 118:53 ICache.scala 118:53]
  wire  _GEN_785 = 5'h6 == index_addr; // @[ICache.scala 118:53 ICache.scala 118:53]
  wire  _GEN_786 = 5'h7 == index_addr; // @[ICache.scala 118:53 ICache.scala 118:53]
  wire  _GEN_787 = 5'h8 == index_addr; // @[ICache.scala 118:53 ICache.scala 118:53]
  wire  _GEN_788 = 5'h9 == index_addr; // @[ICache.scala 118:53 ICache.scala 118:53]
  wire  _GEN_789 = 5'ha == index_addr; // @[ICache.scala 118:53 ICache.scala 118:53]
  wire  _GEN_790 = 5'hb == index_addr; // @[ICache.scala 118:53 ICache.scala 118:53]
  wire  _GEN_791 = 5'hc == index_addr; // @[ICache.scala 118:53 ICache.scala 118:53]
  wire  _GEN_792 = 5'hd == index_addr; // @[ICache.scala 118:53 ICache.scala 118:53]
  wire  _GEN_793 = 5'he == index_addr; // @[ICache.scala 118:53 ICache.scala 118:53]
  wire  _GEN_794 = 5'hf == index_addr; // @[ICache.scala 118:53 ICache.scala 118:53]
  wire  _GEN_795 = 5'h10 == index_addr; // @[ICache.scala 118:53 ICache.scala 118:53]
  wire  _GEN_796 = 5'h11 == index_addr; // @[ICache.scala 118:53 ICache.scala 118:53]
  wire  _GEN_797 = 5'h12 == index_addr; // @[ICache.scala 118:53 ICache.scala 118:53]
  wire  _GEN_798 = 5'h13 == index_addr; // @[ICache.scala 118:53 ICache.scala 118:53]
  wire  _GEN_799 = 5'h14 == index_addr; // @[ICache.scala 118:53 ICache.scala 118:53]
  wire  _GEN_800 = 5'h15 == index_addr; // @[ICache.scala 118:53 ICache.scala 118:53]
  wire  _GEN_801 = 5'h16 == index_addr; // @[ICache.scala 118:53 ICache.scala 118:53]
  wire  _GEN_802 = 5'h17 == index_addr; // @[ICache.scala 118:53 ICache.scala 118:53]
  wire  _GEN_803 = 5'h18 == index_addr; // @[ICache.scala 118:53 ICache.scala 118:53]
  wire  _GEN_804 = 5'h19 == index_addr; // @[ICache.scala 118:53 ICache.scala 118:53]
  wire  _GEN_805 = 5'h1a == index_addr; // @[ICache.scala 118:53 ICache.scala 118:53]
  wire  _GEN_806 = 5'h1b == index_addr; // @[ICache.scala 118:53 ICache.scala 118:53]
  wire  _GEN_807 = 5'h1c == index_addr; // @[ICache.scala 118:53 ICache.scala 118:53]
  wire  _GEN_808 = 5'h1d == index_addr; // @[ICache.scala 118:53 ICache.scala 118:53]
  wire  _GEN_809 = 5'h1e == index_addr; // @[ICache.scala 118:53 ICache.scala 118:53]
  wire  _GEN_810 = 5'h1f == index_addr; // @[ICache.scala 118:53 ICache.scala 118:53]
  wire  _T_11 = state == 2'h3; // @[ICache.scala 119:16]
  wire [4:0] _fence_cnt_T_1 = fence_cnt + 5'h1; // @[ICache.scala 123:83]
  assign io_imem_data = hit2 ? data2 : _data_T; // @[ICache.scala 68:22]
  assign io_imem_ok = (hit | not_en_yet) & state == 2'h0; // @[ICache.scala 82:44]
  assign io_axi_req = state == 2'h1; // @[ICache.scala 102:28]
  assign io_axi_addr = addr & 64'hffffffffffffffc0; // @[ICache.scala 103:27]
  assign io_fence_done = _T_6 & _T_11; // @[ICache.scala 127:57]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 27:20]
      addr <= 64'h0; // @[Reg.scala 27:20]
    end else if (_addr_T) begin // @[Reg.scala 28:19]
      addr <= io_imem_addr; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[ICache.scala 53:26]
      v1_0 <= 1'h0; // @[ICache.scala 53:26]
    end else if (state == 2'h2) begin // @[ICache.scala 117:37]
      if (5'h0 == fence_cnt) begin // @[ICache.scala 117:52]
        v1_0 <= 1'h0; // @[ICache.scala 117:52]
      end else begin
        v1_0 <= _GEN_394;
      end
    end else if (_block1_T) begin // @[ICache.scala 118:37]
      v1_0 <= 5'h0 == index_addr | _GEN_394;
    end else begin
      v1_0 <= _GEN_394;
    end
    if (reset) begin // @[ICache.scala 53:26]
      v1_1 <= 1'h0; // @[ICache.scala 53:26]
    end else if (state == 2'h2) begin // @[ICache.scala 117:37]
      if (5'h1 == fence_cnt) begin // @[ICache.scala 117:52]
        v1_1 <= 1'h0; // @[ICache.scala 117:52]
      end else begin
        v1_1 <= _GEN_395;
      end
    end else if (_block1_T) begin // @[ICache.scala 118:37]
      v1_1 <= 5'h1 == index_addr | _GEN_395;
    end else begin
      v1_1 <= _GEN_395;
    end
    if (reset) begin // @[ICache.scala 53:26]
      v1_2 <= 1'h0; // @[ICache.scala 53:26]
    end else if (state == 2'h2) begin // @[ICache.scala 117:37]
      if (5'h2 == fence_cnt) begin // @[ICache.scala 117:52]
        v1_2 <= 1'h0; // @[ICache.scala 117:52]
      end else begin
        v1_2 <= _GEN_396;
      end
    end else if (_block1_T) begin // @[ICache.scala 118:37]
      v1_2 <= 5'h2 == index_addr | _GEN_396;
    end else begin
      v1_2 <= _GEN_396;
    end
    if (reset) begin // @[ICache.scala 53:26]
      v1_3 <= 1'h0; // @[ICache.scala 53:26]
    end else if (state == 2'h2) begin // @[ICache.scala 117:37]
      if (5'h3 == fence_cnt) begin // @[ICache.scala 117:52]
        v1_3 <= 1'h0; // @[ICache.scala 117:52]
      end else begin
        v1_3 <= _GEN_397;
      end
    end else if (_block1_T) begin // @[ICache.scala 118:37]
      v1_3 <= 5'h3 == index_addr | _GEN_397;
    end else begin
      v1_3 <= _GEN_397;
    end
    if (reset) begin // @[ICache.scala 53:26]
      v1_4 <= 1'h0; // @[ICache.scala 53:26]
    end else if (state == 2'h2) begin // @[ICache.scala 117:37]
      if (5'h4 == fence_cnt) begin // @[ICache.scala 117:52]
        v1_4 <= 1'h0; // @[ICache.scala 117:52]
      end else begin
        v1_4 <= _GEN_398;
      end
    end else if (_block1_T) begin // @[ICache.scala 118:37]
      v1_4 <= 5'h4 == index_addr | _GEN_398;
    end else begin
      v1_4 <= _GEN_398;
    end
    if (reset) begin // @[ICache.scala 53:26]
      v1_5 <= 1'h0; // @[ICache.scala 53:26]
    end else if (state == 2'h2) begin // @[ICache.scala 117:37]
      if (5'h5 == fence_cnt) begin // @[ICache.scala 117:52]
        v1_5 <= 1'h0; // @[ICache.scala 117:52]
      end else begin
        v1_5 <= _GEN_399;
      end
    end else if (_block1_T) begin // @[ICache.scala 118:37]
      v1_5 <= 5'h5 == index_addr | _GEN_399;
    end else begin
      v1_5 <= _GEN_399;
    end
    if (reset) begin // @[ICache.scala 53:26]
      v1_6 <= 1'h0; // @[ICache.scala 53:26]
    end else if (state == 2'h2) begin // @[ICache.scala 117:37]
      if (5'h6 == fence_cnt) begin // @[ICache.scala 117:52]
        v1_6 <= 1'h0; // @[ICache.scala 117:52]
      end else begin
        v1_6 <= _GEN_400;
      end
    end else if (_block1_T) begin // @[ICache.scala 118:37]
      v1_6 <= 5'h6 == index_addr | _GEN_400;
    end else begin
      v1_6 <= _GEN_400;
    end
    if (reset) begin // @[ICache.scala 53:26]
      v1_7 <= 1'h0; // @[ICache.scala 53:26]
    end else if (state == 2'h2) begin // @[ICache.scala 117:37]
      if (5'h7 == fence_cnt) begin // @[ICache.scala 117:52]
        v1_7 <= 1'h0; // @[ICache.scala 117:52]
      end else begin
        v1_7 <= _GEN_401;
      end
    end else if (_block1_T) begin // @[ICache.scala 118:37]
      v1_7 <= 5'h7 == index_addr | _GEN_401;
    end else begin
      v1_7 <= _GEN_401;
    end
    if (reset) begin // @[ICache.scala 53:26]
      v1_8 <= 1'h0; // @[ICache.scala 53:26]
    end else if (state == 2'h2) begin // @[ICache.scala 117:37]
      if (5'h8 == fence_cnt) begin // @[ICache.scala 117:52]
        v1_8 <= 1'h0; // @[ICache.scala 117:52]
      end else begin
        v1_8 <= _GEN_402;
      end
    end else if (_block1_T) begin // @[ICache.scala 118:37]
      v1_8 <= 5'h8 == index_addr | _GEN_402;
    end else begin
      v1_8 <= _GEN_402;
    end
    if (reset) begin // @[ICache.scala 53:26]
      v1_9 <= 1'h0; // @[ICache.scala 53:26]
    end else if (state == 2'h2) begin // @[ICache.scala 117:37]
      if (5'h9 == fence_cnt) begin // @[ICache.scala 117:52]
        v1_9 <= 1'h0; // @[ICache.scala 117:52]
      end else begin
        v1_9 <= _GEN_403;
      end
    end else if (_block1_T) begin // @[ICache.scala 118:37]
      v1_9 <= 5'h9 == index_addr | _GEN_403;
    end else begin
      v1_9 <= _GEN_403;
    end
    if (reset) begin // @[ICache.scala 53:26]
      v1_10 <= 1'h0; // @[ICache.scala 53:26]
    end else if (state == 2'h2) begin // @[ICache.scala 117:37]
      if (5'ha == fence_cnt) begin // @[ICache.scala 117:52]
        v1_10 <= 1'h0; // @[ICache.scala 117:52]
      end else begin
        v1_10 <= _GEN_404;
      end
    end else if (_block1_T) begin // @[ICache.scala 118:37]
      v1_10 <= 5'ha == index_addr | _GEN_404;
    end else begin
      v1_10 <= _GEN_404;
    end
    if (reset) begin // @[ICache.scala 53:26]
      v1_11 <= 1'h0; // @[ICache.scala 53:26]
    end else if (state == 2'h2) begin // @[ICache.scala 117:37]
      if (5'hb == fence_cnt) begin // @[ICache.scala 117:52]
        v1_11 <= 1'h0; // @[ICache.scala 117:52]
      end else begin
        v1_11 <= _GEN_405;
      end
    end else if (_block1_T) begin // @[ICache.scala 118:37]
      v1_11 <= 5'hb == index_addr | _GEN_405;
    end else begin
      v1_11 <= _GEN_405;
    end
    if (reset) begin // @[ICache.scala 53:26]
      v1_12 <= 1'h0; // @[ICache.scala 53:26]
    end else if (state == 2'h2) begin // @[ICache.scala 117:37]
      if (5'hc == fence_cnt) begin // @[ICache.scala 117:52]
        v1_12 <= 1'h0; // @[ICache.scala 117:52]
      end else begin
        v1_12 <= _GEN_406;
      end
    end else if (_block1_T) begin // @[ICache.scala 118:37]
      v1_12 <= 5'hc == index_addr | _GEN_406;
    end else begin
      v1_12 <= _GEN_406;
    end
    if (reset) begin // @[ICache.scala 53:26]
      v1_13 <= 1'h0; // @[ICache.scala 53:26]
    end else if (state == 2'h2) begin // @[ICache.scala 117:37]
      if (5'hd == fence_cnt) begin // @[ICache.scala 117:52]
        v1_13 <= 1'h0; // @[ICache.scala 117:52]
      end else begin
        v1_13 <= _GEN_407;
      end
    end else if (_block1_T) begin // @[ICache.scala 118:37]
      v1_13 <= 5'hd == index_addr | _GEN_407;
    end else begin
      v1_13 <= _GEN_407;
    end
    if (reset) begin // @[ICache.scala 53:26]
      v1_14 <= 1'h0; // @[ICache.scala 53:26]
    end else if (state == 2'h2) begin // @[ICache.scala 117:37]
      if (5'he == fence_cnt) begin // @[ICache.scala 117:52]
        v1_14 <= 1'h0; // @[ICache.scala 117:52]
      end else begin
        v1_14 <= _GEN_408;
      end
    end else if (_block1_T) begin // @[ICache.scala 118:37]
      v1_14 <= 5'he == index_addr | _GEN_408;
    end else begin
      v1_14 <= _GEN_408;
    end
    if (reset) begin // @[ICache.scala 53:26]
      v1_15 <= 1'h0; // @[ICache.scala 53:26]
    end else if (state == 2'h2) begin // @[ICache.scala 117:37]
      if (5'hf == fence_cnt) begin // @[ICache.scala 117:52]
        v1_15 <= 1'h0; // @[ICache.scala 117:52]
      end else begin
        v1_15 <= _GEN_409;
      end
    end else if (_block1_T) begin // @[ICache.scala 118:37]
      v1_15 <= 5'hf == index_addr | _GEN_409;
    end else begin
      v1_15 <= _GEN_409;
    end
    if (reset) begin // @[ICache.scala 53:26]
      v1_16 <= 1'h0; // @[ICache.scala 53:26]
    end else if (state == 2'h2) begin // @[ICache.scala 117:37]
      if (5'h10 == fence_cnt) begin // @[ICache.scala 117:52]
        v1_16 <= 1'h0; // @[ICache.scala 117:52]
      end else begin
        v1_16 <= _GEN_410;
      end
    end else if (_block1_T) begin // @[ICache.scala 118:37]
      v1_16 <= 5'h10 == index_addr | _GEN_410;
    end else begin
      v1_16 <= _GEN_410;
    end
    if (reset) begin // @[ICache.scala 53:26]
      v1_17 <= 1'h0; // @[ICache.scala 53:26]
    end else if (state == 2'h2) begin // @[ICache.scala 117:37]
      if (5'h11 == fence_cnt) begin // @[ICache.scala 117:52]
        v1_17 <= 1'h0; // @[ICache.scala 117:52]
      end else begin
        v1_17 <= _GEN_411;
      end
    end else if (_block1_T) begin // @[ICache.scala 118:37]
      v1_17 <= 5'h11 == index_addr | _GEN_411;
    end else begin
      v1_17 <= _GEN_411;
    end
    if (reset) begin // @[ICache.scala 53:26]
      v1_18 <= 1'h0; // @[ICache.scala 53:26]
    end else if (state == 2'h2) begin // @[ICache.scala 117:37]
      if (5'h12 == fence_cnt) begin // @[ICache.scala 117:52]
        v1_18 <= 1'h0; // @[ICache.scala 117:52]
      end else begin
        v1_18 <= _GEN_412;
      end
    end else if (_block1_T) begin // @[ICache.scala 118:37]
      v1_18 <= 5'h12 == index_addr | _GEN_412;
    end else begin
      v1_18 <= _GEN_412;
    end
    if (reset) begin // @[ICache.scala 53:26]
      v1_19 <= 1'h0; // @[ICache.scala 53:26]
    end else if (state == 2'h2) begin // @[ICache.scala 117:37]
      if (5'h13 == fence_cnt) begin // @[ICache.scala 117:52]
        v1_19 <= 1'h0; // @[ICache.scala 117:52]
      end else begin
        v1_19 <= _GEN_413;
      end
    end else if (_block1_T) begin // @[ICache.scala 118:37]
      v1_19 <= 5'h13 == index_addr | _GEN_413;
    end else begin
      v1_19 <= _GEN_413;
    end
    if (reset) begin // @[ICache.scala 53:26]
      v1_20 <= 1'h0; // @[ICache.scala 53:26]
    end else if (state == 2'h2) begin // @[ICache.scala 117:37]
      if (5'h14 == fence_cnt) begin // @[ICache.scala 117:52]
        v1_20 <= 1'h0; // @[ICache.scala 117:52]
      end else begin
        v1_20 <= _GEN_414;
      end
    end else if (_block1_T) begin // @[ICache.scala 118:37]
      v1_20 <= 5'h14 == index_addr | _GEN_414;
    end else begin
      v1_20 <= _GEN_414;
    end
    if (reset) begin // @[ICache.scala 53:26]
      v1_21 <= 1'h0; // @[ICache.scala 53:26]
    end else if (state == 2'h2) begin // @[ICache.scala 117:37]
      if (5'h15 == fence_cnt) begin // @[ICache.scala 117:52]
        v1_21 <= 1'h0; // @[ICache.scala 117:52]
      end else begin
        v1_21 <= _GEN_415;
      end
    end else if (_block1_T) begin // @[ICache.scala 118:37]
      v1_21 <= 5'h15 == index_addr | _GEN_415;
    end else begin
      v1_21 <= _GEN_415;
    end
    if (reset) begin // @[ICache.scala 53:26]
      v1_22 <= 1'h0; // @[ICache.scala 53:26]
    end else if (state == 2'h2) begin // @[ICache.scala 117:37]
      if (5'h16 == fence_cnt) begin // @[ICache.scala 117:52]
        v1_22 <= 1'h0; // @[ICache.scala 117:52]
      end else begin
        v1_22 <= _GEN_416;
      end
    end else if (_block1_T) begin // @[ICache.scala 118:37]
      v1_22 <= 5'h16 == index_addr | _GEN_416;
    end else begin
      v1_22 <= _GEN_416;
    end
    if (reset) begin // @[ICache.scala 53:26]
      v1_23 <= 1'h0; // @[ICache.scala 53:26]
    end else if (state == 2'h2) begin // @[ICache.scala 117:37]
      if (5'h17 == fence_cnt) begin // @[ICache.scala 117:52]
        v1_23 <= 1'h0; // @[ICache.scala 117:52]
      end else begin
        v1_23 <= _GEN_417;
      end
    end else if (_block1_T) begin // @[ICache.scala 118:37]
      v1_23 <= 5'h17 == index_addr | _GEN_417;
    end else begin
      v1_23 <= _GEN_417;
    end
    if (reset) begin // @[ICache.scala 53:26]
      v1_24 <= 1'h0; // @[ICache.scala 53:26]
    end else if (state == 2'h2) begin // @[ICache.scala 117:37]
      if (5'h18 == fence_cnt) begin // @[ICache.scala 117:52]
        v1_24 <= 1'h0; // @[ICache.scala 117:52]
      end else begin
        v1_24 <= _GEN_418;
      end
    end else if (_block1_T) begin // @[ICache.scala 118:37]
      v1_24 <= 5'h18 == index_addr | _GEN_418;
    end else begin
      v1_24 <= _GEN_418;
    end
    if (reset) begin // @[ICache.scala 53:26]
      v1_25 <= 1'h0; // @[ICache.scala 53:26]
    end else if (state == 2'h2) begin // @[ICache.scala 117:37]
      if (5'h19 == fence_cnt) begin // @[ICache.scala 117:52]
        v1_25 <= 1'h0; // @[ICache.scala 117:52]
      end else begin
        v1_25 <= _GEN_419;
      end
    end else if (_block1_T) begin // @[ICache.scala 118:37]
      v1_25 <= 5'h19 == index_addr | _GEN_419;
    end else begin
      v1_25 <= _GEN_419;
    end
    if (reset) begin // @[ICache.scala 53:26]
      v1_26 <= 1'h0; // @[ICache.scala 53:26]
    end else if (state == 2'h2) begin // @[ICache.scala 117:37]
      if (5'h1a == fence_cnt) begin // @[ICache.scala 117:52]
        v1_26 <= 1'h0; // @[ICache.scala 117:52]
      end else begin
        v1_26 <= _GEN_420;
      end
    end else if (_block1_T) begin // @[ICache.scala 118:37]
      v1_26 <= 5'h1a == index_addr | _GEN_420;
    end else begin
      v1_26 <= _GEN_420;
    end
    if (reset) begin // @[ICache.scala 53:26]
      v1_27 <= 1'h0; // @[ICache.scala 53:26]
    end else if (state == 2'h2) begin // @[ICache.scala 117:37]
      if (5'h1b == fence_cnt) begin // @[ICache.scala 117:52]
        v1_27 <= 1'h0; // @[ICache.scala 117:52]
      end else begin
        v1_27 <= _GEN_421;
      end
    end else if (_block1_T) begin // @[ICache.scala 118:37]
      v1_27 <= 5'h1b == index_addr | _GEN_421;
    end else begin
      v1_27 <= _GEN_421;
    end
    if (reset) begin // @[ICache.scala 53:26]
      v1_28 <= 1'h0; // @[ICache.scala 53:26]
    end else if (state == 2'h2) begin // @[ICache.scala 117:37]
      if (5'h1c == fence_cnt) begin // @[ICache.scala 117:52]
        v1_28 <= 1'h0; // @[ICache.scala 117:52]
      end else begin
        v1_28 <= _GEN_422;
      end
    end else if (_block1_T) begin // @[ICache.scala 118:37]
      v1_28 <= 5'h1c == index_addr | _GEN_422;
    end else begin
      v1_28 <= _GEN_422;
    end
    if (reset) begin // @[ICache.scala 53:26]
      v1_29 <= 1'h0; // @[ICache.scala 53:26]
    end else if (state == 2'h2) begin // @[ICache.scala 117:37]
      if (5'h1d == fence_cnt) begin // @[ICache.scala 117:52]
        v1_29 <= 1'h0; // @[ICache.scala 117:52]
      end else begin
        v1_29 <= _GEN_423;
      end
    end else if (_block1_T) begin // @[ICache.scala 118:37]
      v1_29 <= 5'h1d == index_addr | _GEN_423;
    end else begin
      v1_29 <= _GEN_423;
    end
    if (reset) begin // @[ICache.scala 53:26]
      v1_30 <= 1'h0; // @[ICache.scala 53:26]
    end else if (state == 2'h2) begin // @[ICache.scala 117:37]
      if (5'h1e == fence_cnt) begin // @[ICache.scala 117:52]
        v1_30 <= 1'h0; // @[ICache.scala 117:52]
      end else begin
        v1_30 <= _GEN_424;
      end
    end else if (_block1_T) begin // @[ICache.scala 118:37]
      v1_30 <= 5'h1e == index_addr | _GEN_424;
    end else begin
      v1_30 <= _GEN_424;
    end
    if (reset) begin // @[ICache.scala 53:26]
      v1_31 <= 1'h0; // @[ICache.scala 53:26]
    end else if (state == 2'h2) begin // @[ICache.scala 117:37]
      if (5'h1f == fence_cnt) begin // @[ICache.scala 117:52]
        v1_31 <= 1'h0; // @[ICache.scala 117:52]
      end else begin
        v1_31 <= _GEN_425;
      end
    end else if (_block1_T) begin // @[ICache.scala 118:37]
      v1_31 <= 5'h1f == index_addr | _GEN_425;
    end else begin
      v1_31 <= _GEN_425;
    end
    if (reset) begin // @[ICache.scala 54:26]
      age1_0 <= 1'h0; // @[ICache.scala 54:26]
    end else if (5'h0 == index_addr) begin // @[ICache.scala 71:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 71:28]
        age1_0 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 71:28]
        age1_0 <= age1_31; // @[ICache.scala 71:28]
      end else begin
        age1_0 <= _GEN_223;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      age1_1 <= 1'h0; // @[ICache.scala 54:26]
    end else if (5'h1 == index_addr) begin // @[ICache.scala 71:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 71:28]
        age1_1 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 71:28]
        age1_1 <= age1_31; // @[ICache.scala 71:28]
      end else begin
        age1_1 <= _GEN_223;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      age1_2 <= 1'h0; // @[ICache.scala 54:26]
    end else if (5'h2 == index_addr) begin // @[ICache.scala 71:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 71:28]
        age1_2 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 71:28]
        age1_2 <= age1_31; // @[ICache.scala 71:28]
      end else begin
        age1_2 <= _GEN_223;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      age1_3 <= 1'h0; // @[ICache.scala 54:26]
    end else if (5'h3 == index_addr) begin // @[ICache.scala 71:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 71:28]
        age1_3 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 71:28]
        age1_3 <= age1_31; // @[ICache.scala 71:28]
      end else begin
        age1_3 <= _GEN_223;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      age1_4 <= 1'h0; // @[ICache.scala 54:26]
    end else if (5'h4 == index_addr) begin // @[ICache.scala 71:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 71:28]
        age1_4 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 71:28]
        age1_4 <= age1_31; // @[ICache.scala 71:28]
      end else begin
        age1_4 <= _GEN_223;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      age1_5 <= 1'h0; // @[ICache.scala 54:26]
    end else if (5'h5 == index_addr) begin // @[ICache.scala 71:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 71:28]
        age1_5 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 71:28]
        age1_5 <= age1_31; // @[ICache.scala 71:28]
      end else begin
        age1_5 <= _GEN_223;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      age1_6 <= 1'h0; // @[ICache.scala 54:26]
    end else if (5'h6 == index_addr) begin // @[ICache.scala 71:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 71:28]
        age1_6 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 71:28]
        age1_6 <= age1_31; // @[ICache.scala 71:28]
      end else begin
        age1_6 <= _GEN_223;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      age1_7 <= 1'h0; // @[ICache.scala 54:26]
    end else if (5'h7 == index_addr) begin // @[ICache.scala 71:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 71:28]
        age1_7 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 71:28]
        age1_7 <= age1_31; // @[ICache.scala 71:28]
      end else begin
        age1_7 <= _GEN_223;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      age1_8 <= 1'h0; // @[ICache.scala 54:26]
    end else if (5'h8 == index_addr) begin // @[ICache.scala 71:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 71:28]
        age1_8 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 71:28]
        age1_8 <= age1_31; // @[ICache.scala 71:28]
      end else begin
        age1_8 <= _GEN_223;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      age1_9 <= 1'h0; // @[ICache.scala 54:26]
    end else if (5'h9 == index_addr) begin // @[ICache.scala 71:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 71:28]
        age1_9 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 71:28]
        age1_9 <= age1_31; // @[ICache.scala 71:28]
      end else begin
        age1_9 <= _GEN_223;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      age1_10 <= 1'h0; // @[ICache.scala 54:26]
    end else if (5'ha == index_addr) begin // @[ICache.scala 71:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 71:28]
        age1_10 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 71:28]
        age1_10 <= age1_31; // @[ICache.scala 71:28]
      end else begin
        age1_10 <= _GEN_223;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      age1_11 <= 1'h0; // @[ICache.scala 54:26]
    end else if (5'hb == index_addr) begin // @[ICache.scala 71:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 71:28]
        age1_11 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 71:28]
        age1_11 <= age1_31; // @[ICache.scala 71:28]
      end else begin
        age1_11 <= _GEN_223;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      age1_12 <= 1'h0; // @[ICache.scala 54:26]
    end else if (5'hc == index_addr) begin // @[ICache.scala 71:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 71:28]
        age1_12 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 71:28]
        age1_12 <= age1_31; // @[ICache.scala 71:28]
      end else begin
        age1_12 <= _GEN_223;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      age1_13 <= 1'h0; // @[ICache.scala 54:26]
    end else if (5'hd == index_addr) begin // @[ICache.scala 71:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 71:28]
        age1_13 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 71:28]
        age1_13 <= age1_31; // @[ICache.scala 71:28]
      end else begin
        age1_13 <= _GEN_223;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      age1_14 <= 1'h0; // @[ICache.scala 54:26]
    end else if (5'he == index_addr) begin // @[ICache.scala 71:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 71:28]
        age1_14 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 71:28]
        age1_14 <= age1_31; // @[ICache.scala 71:28]
      end else begin
        age1_14 <= _GEN_223;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      age1_15 <= 1'h0; // @[ICache.scala 54:26]
    end else if (5'hf == index_addr) begin // @[ICache.scala 71:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 71:28]
        age1_15 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 71:28]
        age1_15 <= age1_31; // @[ICache.scala 71:28]
      end else begin
        age1_15 <= _GEN_223;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      age1_16 <= 1'h0; // @[ICache.scala 54:26]
    end else if (5'h10 == index_addr) begin // @[ICache.scala 71:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 71:28]
        age1_16 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 71:28]
        age1_16 <= age1_31; // @[ICache.scala 71:28]
      end else begin
        age1_16 <= _GEN_223;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      age1_17 <= 1'h0; // @[ICache.scala 54:26]
    end else if (5'h11 == index_addr) begin // @[ICache.scala 71:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 71:28]
        age1_17 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 71:28]
        age1_17 <= age1_31; // @[ICache.scala 71:28]
      end else begin
        age1_17 <= _GEN_223;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      age1_18 <= 1'h0; // @[ICache.scala 54:26]
    end else if (5'h12 == index_addr) begin // @[ICache.scala 71:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 71:28]
        age1_18 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 71:28]
        age1_18 <= age1_31; // @[ICache.scala 71:28]
      end else begin
        age1_18 <= _GEN_223;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      age1_19 <= 1'h0; // @[ICache.scala 54:26]
    end else if (5'h13 == index_addr) begin // @[ICache.scala 71:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 71:28]
        age1_19 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 71:28]
        age1_19 <= age1_31; // @[ICache.scala 71:28]
      end else begin
        age1_19 <= _GEN_223;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      age1_20 <= 1'h0; // @[ICache.scala 54:26]
    end else if (5'h14 == index_addr) begin // @[ICache.scala 71:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 71:28]
        age1_20 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 71:28]
        age1_20 <= age1_31; // @[ICache.scala 71:28]
      end else begin
        age1_20 <= _GEN_223;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      age1_21 <= 1'h0; // @[ICache.scala 54:26]
    end else if (5'h15 == index_addr) begin // @[ICache.scala 71:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 71:28]
        age1_21 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 71:28]
        age1_21 <= age1_31; // @[ICache.scala 71:28]
      end else begin
        age1_21 <= _GEN_223;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      age1_22 <= 1'h0; // @[ICache.scala 54:26]
    end else if (5'h16 == index_addr) begin // @[ICache.scala 71:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 71:28]
        age1_22 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 71:28]
        age1_22 <= age1_31; // @[ICache.scala 71:28]
      end else begin
        age1_22 <= _GEN_223;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      age1_23 <= 1'h0; // @[ICache.scala 54:26]
    end else if (5'h17 == index_addr) begin // @[ICache.scala 71:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 71:28]
        age1_23 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 71:28]
        age1_23 <= age1_31; // @[ICache.scala 71:28]
      end else begin
        age1_23 <= _GEN_223;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      age1_24 <= 1'h0; // @[ICache.scala 54:26]
    end else if (5'h18 == index_addr) begin // @[ICache.scala 71:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 71:28]
        age1_24 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 71:28]
        age1_24 <= age1_31; // @[ICache.scala 71:28]
      end else begin
        age1_24 <= _GEN_223;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      age1_25 <= 1'h0; // @[ICache.scala 54:26]
    end else if (5'h19 == index_addr) begin // @[ICache.scala 71:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 71:28]
        age1_25 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 71:28]
        age1_25 <= age1_31; // @[ICache.scala 71:28]
      end else begin
        age1_25 <= _GEN_223;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      age1_26 <= 1'h0; // @[ICache.scala 54:26]
    end else if (5'h1a == index_addr) begin // @[ICache.scala 71:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 71:28]
        age1_26 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 71:28]
        age1_26 <= age1_31; // @[ICache.scala 71:28]
      end else begin
        age1_26 <= _GEN_223;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      age1_27 <= 1'h0; // @[ICache.scala 54:26]
    end else if (5'h1b == index_addr) begin // @[ICache.scala 71:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 71:28]
        age1_27 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 71:28]
        age1_27 <= age1_31; // @[ICache.scala 71:28]
      end else begin
        age1_27 <= _GEN_223;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      age1_28 <= 1'h0; // @[ICache.scala 54:26]
    end else if (5'h1c == index_addr) begin // @[ICache.scala 71:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 71:28]
        age1_28 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 71:28]
        age1_28 <= age1_31; // @[ICache.scala 71:28]
      end else begin
        age1_28 <= _GEN_223;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      age1_29 <= 1'h0; // @[ICache.scala 54:26]
    end else if (5'h1d == index_addr) begin // @[ICache.scala 71:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 71:28]
        age1_29 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 71:28]
        age1_29 <= age1_31; // @[ICache.scala 71:28]
      end else begin
        age1_29 <= _GEN_223;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      age1_30 <= 1'h0; // @[ICache.scala 54:26]
    end else if (5'h1e == index_addr) begin // @[ICache.scala 71:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 71:28]
        age1_30 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 71:28]
        age1_30 <= age1_31; // @[ICache.scala 71:28]
      end else begin
        age1_30 <= _GEN_223;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      age1_31 <= 1'h0; // @[ICache.scala 54:26]
    end else if (5'h1f == index_addr) begin // @[ICache.scala 71:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 71:28]
        age1_31 <= hit1;
      end else if (!(5'h1f == index_addr)) begin // @[ICache.scala 71:28]
        age1_31 <= _GEN_223;
      end
    end
    if (reset) begin // @[ICache.scala 55:26]
      tag1_0 <= 53'h0; // @[ICache.scala 55:26]
    end else if (5'h0 == index_addr) begin // @[ICache.scala 111:26]
      if (_block1_T) begin // @[ICache.scala 111:32]
        tag1_0 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 62:28]
        tag1_0 <= tag1_31; // @[ICache.scala 62:28]
      end else begin
        tag1_0 <= _GEN_31;
      end
    end
    if (reset) begin // @[ICache.scala 55:26]
      tag1_1 <= 53'h0; // @[ICache.scala 55:26]
    end else if (5'h1 == index_addr) begin // @[ICache.scala 111:26]
      if (_block1_T) begin // @[ICache.scala 111:32]
        tag1_1 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 62:28]
        tag1_1 <= tag1_31; // @[ICache.scala 62:28]
      end else begin
        tag1_1 <= _GEN_31;
      end
    end
    if (reset) begin // @[ICache.scala 55:26]
      tag1_2 <= 53'h0; // @[ICache.scala 55:26]
    end else if (5'h2 == index_addr) begin // @[ICache.scala 111:26]
      if (_block1_T) begin // @[ICache.scala 111:32]
        tag1_2 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 62:28]
        tag1_2 <= tag1_31; // @[ICache.scala 62:28]
      end else begin
        tag1_2 <= _GEN_31;
      end
    end
    if (reset) begin // @[ICache.scala 55:26]
      tag1_3 <= 53'h0; // @[ICache.scala 55:26]
    end else if (5'h3 == index_addr) begin // @[ICache.scala 111:26]
      if (_block1_T) begin // @[ICache.scala 111:32]
        tag1_3 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 62:28]
        tag1_3 <= tag1_31; // @[ICache.scala 62:28]
      end else begin
        tag1_3 <= _GEN_31;
      end
    end
    if (reset) begin // @[ICache.scala 55:26]
      tag1_4 <= 53'h0; // @[ICache.scala 55:26]
    end else if (5'h4 == index_addr) begin // @[ICache.scala 111:26]
      if (_block1_T) begin // @[ICache.scala 111:32]
        tag1_4 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 62:28]
        tag1_4 <= tag1_31; // @[ICache.scala 62:28]
      end else begin
        tag1_4 <= _GEN_31;
      end
    end
    if (reset) begin // @[ICache.scala 55:26]
      tag1_5 <= 53'h0; // @[ICache.scala 55:26]
    end else if (5'h5 == index_addr) begin // @[ICache.scala 111:26]
      if (_block1_T) begin // @[ICache.scala 111:32]
        tag1_5 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 62:28]
        tag1_5 <= tag1_31; // @[ICache.scala 62:28]
      end else begin
        tag1_5 <= _GEN_31;
      end
    end
    if (reset) begin // @[ICache.scala 55:26]
      tag1_6 <= 53'h0; // @[ICache.scala 55:26]
    end else if (5'h6 == index_addr) begin // @[ICache.scala 111:26]
      if (_block1_T) begin // @[ICache.scala 111:32]
        tag1_6 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 62:28]
        tag1_6 <= tag1_31; // @[ICache.scala 62:28]
      end else begin
        tag1_6 <= _GEN_31;
      end
    end
    if (reset) begin // @[ICache.scala 55:26]
      tag1_7 <= 53'h0; // @[ICache.scala 55:26]
    end else if (5'h7 == index_addr) begin // @[ICache.scala 111:26]
      if (_block1_T) begin // @[ICache.scala 111:32]
        tag1_7 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 62:28]
        tag1_7 <= tag1_31; // @[ICache.scala 62:28]
      end else begin
        tag1_7 <= _GEN_31;
      end
    end
    if (reset) begin // @[ICache.scala 55:26]
      tag1_8 <= 53'h0; // @[ICache.scala 55:26]
    end else if (5'h8 == index_addr) begin // @[ICache.scala 111:26]
      if (_block1_T) begin // @[ICache.scala 111:32]
        tag1_8 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 62:28]
        tag1_8 <= tag1_31; // @[ICache.scala 62:28]
      end else begin
        tag1_8 <= _GEN_31;
      end
    end
    if (reset) begin // @[ICache.scala 55:26]
      tag1_9 <= 53'h0; // @[ICache.scala 55:26]
    end else if (5'h9 == index_addr) begin // @[ICache.scala 111:26]
      if (_block1_T) begin // @[ICache.scala 111:32]
        tag1_9 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 62:28]
        tag1_9 <= tag1_31; // @[ICache.scala 62:28]
      end else begin
        tag1_9 <= _GEN_31;
      end
    end
    if (reset) begin // @[ICache.scala 55:26]
      tag1_10 <= 53'h0; // @[ICache.scala 55:26]
    end else if (5'ha == index_addr) begin // @[ICache.scala 111:26]
      if (_block1_T) begin // @[ICache.scala 111:32]
        tag1_10 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 62:28]
        tag1_10 <= tag1_31; // @[ICache.scala 62:28]
      end else begin
        tag1_10 <= _GEN_31;
      end
    end
    if (reset) begin // @[ICache.scala 55:26]
      tag1_11 <= 53'h0; // @[ICache.scala 55:26]
    end else if (5'hb == index_addr) begin // @[ICache.scala 111:26]
      if (_block1_T) begin // @[ICache.scala 111:32]
        tag1_11 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 62:28]
        tag1_11 <= tag1_31; // @[ICache.scala 62:28]
      end else begin
        tag1_11 <= _GEN_31;
      end
    end
    if (reset) begin // @[ICache.scala 55:26]
      tag1_12 <= 53'h0; // @[ICache.scala 55:26]
    end else if (5'hc == index_addr) begin // @[ICache.scala 111:26]
      if (_block1_T) begin // @[ICache.scala 111:32]
        tag1_12 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 62:28]
        tag1_12 <= tag1_31; // @[ICache.scala 62:28]
      end else begin
        tag1_12 <= _GEN_31;
      end
    end
    if (reset) begin // @[ICache.scala 55:26]
      tag1_13 <= 53'h0; // @[ICache.scala 55:26]
    end else if (5'hd == index_addr) begin // @[ICache.scala 111:26]
      if (_block1_T) begin // @[ICache.scala 111:32]
        tag1_13 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 62:28]
        tag1_13 <= tag1_31; // @[ICache.scala 62:28]
      end else begin
        tag1_13 <= _GEN_31;
      end
    end
    if (reset) begin // @[ICache.scala 55:26]
      tag1_14 <= 53'h0; // @[ICache.scala 55:26]
    end else if (5'he == index_addr) begin // @[ICache.scala 111:26]
      if (_block1_T) begin // @[ICache.scala 111:32]
        tag1_14 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 62:28]
        tag1_14 <= tag1_31; // @[ICache.scala 62:28]
      end else begin
        tag1_14 <= _GEN_31;
      end
    end
    if (reset) begin // @[ICache.scala 55:26]
      tag1_15 <= 53'h0; // @[ICache.scala 55:26]
    end else if (5'hf == index_addr) begin // @[ICache.scala 111:26]
      if (_block1_T) begin // @[ICache.scala 111:32]
        tag1_15 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 62:28]
        tag1_15 <= tag1_31; // @[ICache.scala 62:28]
      end else begin
        tag1_15 <= _GEN_31;
      end
    end
    if (reset) begin // @[ICache.scala 55:26]
      tag1_16 <= 53'h0; // @[ICache.scala 55:26]
    end else if (5'h10 == index_addr) begin // @[ICache.scala 111:26]
      if (_block1_T) begin // @[ICache.scala 111:32]
        tag1_16 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 62:28]
        tag1_16 <= tag1_31; // @[ICache.scala 62:28]
      end else begin
        tag1_16 <= _GEN_31;
      end
    end
    if (reset) begin // @[ICache.scala 55:26]
      tag1_17 <= 53'h0; // @[ICache.scala 55:26]
    end else if (5'h11 == index_addr) begin // @[ICache.scala 111:26]
      if (_block1_T) begin // @[ICache.scala 111:32]
        tag1_17 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 62:28]
        tag1_17 <= tag1_31; // @[ICache.scala 62:28]
      end else begin
        tag1_17 <= _GEN_31;
      end
    end
    if (reset) begin // @[ICache.scala 55:26]
      tag1_18 <= 53'h0; // @[ICache.scala 55:26]
    end else if (5'h12 == index_addr) begin // @[ICache.scala 111:26]
      if (_block1_T) begin // @[ICache.scala 111:32]
        tag1_18 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 62:28]
        tag1_18 <= tag1_31; // @[ICache.scala 62:28]
      end else begin
        tag1_18 <= _GEN_31;
      end
    end
    if (reset) begin // @[ICache.scala 55:26]
      tag1_19 <= 53'h0; // @[ICache.scala 55:26]
    end else if (5'h13 == index_addr) begin // @[ICache.scala 111:26]
      if (_block1_T) begin // @[ICache.scala 111:32]
        tag1_19 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 62:28]
        tag1_19 <= tag1_31; // @[ICache.scala 62:28]
      end else begin
        tag1_19 <= _GEN_31;
      end
    end
    if (reset) begin // @[ICache.scala 55:26]
      tag1_20 <= 53'h0; // @[ICache.scala 55:26]
    end else if (5'h14 == index_addr) begin // @[ICache.scala 111:26]
      if (_block1_T) begin // @[ICache.scala 111:32]
        tag1_20 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 62:28]
        tag1_20 <= tag1_31; // @[ICache.scala 62:28]
      end else begin
        tag1_20 <= _GEN_31;
      end
    end
    if (reset) begin // @[ICache.scala 55:26]
      tag1_21 <= 53'h0; // @[ICache.scala 55:26]
    end else if (5'h15 == index_addr) begin // @[ICache.scala 111:26]
      if (_block1_T) begin // @[ICache.scala 111:32]
        tag1_21 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 62:28]
        tag1_21 <= tag1_31; // @[ICache.scala 62:28]
      end else begin
        tag1_21 <= _GEN_31;
      end
    end
    if (reset) begin // @[ICache.scala 55:26]
      tag1_22 <= 53'h0; // @[ICache.scala 55:26]
    end else if (5'h16 == index_addr) begin // @[ICache.scala 111:26]
      if (_block1_T) begin // @[ICache.scala 111:32]
        tag1_22 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 62:28]
        tag1_22 <= tag1_31; // @[ICache.scala 62:28]
      end else begin
        tag1_22 <= _GEN_31;
      end
    end
    if (reset) begin // @[ICache.scala 55:26]
      tag1_23 <= 53'h0; // @[ICache.scala 55:26]
    end else if (5'h17 == index_addr) begin // @[ICache.scala 111:26]
      if (_block1_T) begin // @[ICache.scala 111:32]
        tag1_23 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 62:28]
        tag1_23 <= tag1_31; // @[ICache.scala 62:28]
      end else begin
        tag1_23 <= _GEN_31;
      end
    end
    if (reset) begin // @[ICache.scala 55:26]
      tag1_24 <= 53'h0; // @[ICache.scala 55:26]
    end else if (5'h18 == index_addr) begin // @[ICache.scala 111:26]
      if (_block1_T) begin // @[ICache.scala 111:32]
        tag1_24 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 62:28]
        tag1_24 <= tag1_31; // @[ICache.scala 62:28]
      end else begin
        tag1_24 <= _GEN_31;
      end
    end
    if (reset) begin // @[ICache.scala 55:26]
      tag1_25 <= 53'h0; // @[ICache.scala 55:26]
    end else if (5'h19 == index_addr) begin // @[ICache.scala 111:26]
      if (_block1_T) begin // @[ICache.scala 111:32]
        tag1_25 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 62:28]
        tag1_25 <= tag1_31; // @[ICache.scala 62:28]
      end else begin
        tag1_25 <= _GEN_31;
      end
    end
    if (reset) begin // @[ICache.scala 55:26]
      tag1_26 <= 53'h0; // @[ICache.scala 55:26]
    end else if (5'h1a == index_addr) begin // @[ICache.scala 111:26]
      if (_block1_T) begin // @[ICache.scala 111:32]
        tag1_26 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 62:28]
        tag1_26 <= tag1_31; // @[ICache.scala 62:28]
      end else begin
        tag1_26 <= _GEN_31;
      end
    end
    if (reset) begin // @[ICache.scala 55:26]
      tag1_27 <= 53'h0; // @[ICache.scala 55:26]
    end else if (5'h1b == index_addr) begin // @[ICache.scala 111:26]
      if (_block1_T) begin // @[ICache.scala 111:32]
        tag1_27 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 62:28]
        tag1_27 <= tag1_31; // @[ICache.scala 62:28]
      end else begin
        tag1_27 <= _GEN_31;
      end
    end
    if (reset) begin // @[ICache.scala 55:26]
      tag1_28 <= 53'h0; // @[ICache.scala 55:26]
    end else if (5'h1c == index_addr) begin // @[ICache.scala 111:26]
      if (_block1_T) begin // @[ICache.scala 111:32]
        tag1_28 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 62:28]
        tag1_28 <= tag1_31; // @[ICache.scala 62:28]
      end else begin
        tag1_28 <= _GEN_31;
      end
    end
    if (reset) begin // @[ICache.scala 55:26]
      tag1_29 <= 53'h0; // @[ICache.scala 55:26]
    end else if (5'h1d == index_addr) begin // @[ICache.scala 111:26]
      if (_block1_T) begin // @[ICache.scala 111:32]
        tag1_29 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 62:28]
        tag1_29 <= tag1_31; // @[ICache.scala 62:28]
      end else begin
        tag1_29 <= _GEN_31;
      end
    end
    if (reset) begin // @[ICache.scala 55:26]
      tag1_30 <= 53'h0; // @[ICache.scala 55:26]
    end else if (5'h1e == index_addr) begin // @[ICache.scala 111:26]
      if (_block1_T) begin // @[ICache.scala 111:32]
        tag1_30 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 62:28]
        tag1_30 <= tag1_31; // @[ICache.scala 62:28]
      end else begin
        tag1_30 <= _GEN_31;
      end
    end
    if (reset) begin // @[ICache.scala 55:26]
      tag1_31 <= 53'h0; // @[ICache.scala 55:26]
    end else if (5'h1f == index_addr) begin // @[ICache.scala 111:26]
      if (_block1_T) begin // @[ICache.scala 111:32]
        tag1_31 <= tag_addr;
      end else if (!(5'h1f == index_addr)) begin // @[ICache.scala 62:28]
        tag1_31 <= _GEN_31;
      end
    end
    if (reset) begin // @[ICache.scala 56:26]
      block1_0 <= 512'h0; // @[ICache.scala 56:26]
    end else if (5'h0 == index_addr) begin // @[ICache.scala 110:26]
      if (update & updateway1) begin // @[ICache.scala 110:32]
        block1_0 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 64:39]
        block1_0 <= block1_31; // @[ICache.scala 64:39]
      end else begin
        block1_0 <= _GEN_159;
      end
    end
    if (reset) begin // @[ICache.scala 56:26]
      block1_1 <= 512'h0; // @[ICache.scala 56:26]
    end else if (5'h1 == index_addr) begin // @[ICache.scala 110:26]
      if (update & updateway1) begin // @[ICache.scala 110:32]
        block1_1 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 64:39]
        block1_1 <= block1_31; // @[ICache.scala 64:39]
      end else begin
        block1_1 <= _GEN_159;
      end
    end
    if (reset) begin // @[ICache.scala 56:26]
      block1_2 <= 512'h0; // @[ICache.scala 56:26]
    end else if (5'h2 == index_addr) begin // @[ICache.scala 110:26]
      if (update & updateway1) begin // @[ICache.scala 110:32]
        block1_2 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 64:39]
        block1_2 <= block1_31; // @[ICache.scala 64:39]
      end else begin
        block1_2 <= _GEN_159;
      end
    end
    if (reset) begin // @[ICache.scala 56:26]
      block1_3 <= 512'h0; // @[ICache.scala 56:26]
    end else if (5'h3 == index_addr) begin // @[ICache.scala 110:26]
      if (update & updateway1) begin // @[ICache.scala 110:32]
        block1_3 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 64:39]
        block1_3 <= block1_31; // @[ICache.scala 64:39]
      end else begin
        block1_3 <= _GEN_159;
      end
    end
    if (reset) begin // @[ICache.scala 56:26]
      block1_4 <= 512'h0; // @[ICache.scala 56:26]
    end else if (5'h4 == index_addr) begin // @[ICache.scala 110:26]
      if (update & updateway1) begin // @[ICache.scala 110:32]
        block1_4 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 64:39]
        block1_4 <= block1_31; // @[ICache.scala 64:39]
      end else begin
        block1_4 <= _GEN_159;
      end
    end
    if (reset) begin // @[ICache.scala 56:26]
      block1_5 <= 512'h0; // @[ICache.scala 56:26]
    end else if (5'h5 == index_addr) begin // @[ICache.scala 110:26]
      if (update & updateway1) begin // @[ICache.scala 110:32]
        block1_5 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 64:39]
        block1_5 <= block1_31; // @[ICache.scala 64:39]
      end else begin
        block1_5 <= _GEN_159;
      end
    end
    if (reset) begin // @[ICache.scala 56:26]
      block1_6 <= 512'h0; // @[ICache.scala 56:26]
    end else if (5'h6 == index_addr) begin // @[ICache.scala 110:26]
      if (update & updateway1) begin // @[ICache.scala 110:32]
        block1_6 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 64:39]
        block1_6 <= block1_31; // @[ICache.scala 64:39]
      end else begin
        block1_6 <= _GEN_159;
      end
    end
    if (reset) begin // @[ICache.scala 56:26]
      block1_7 <= 512'h0; // @[ICache.scala 56:26]
    end else if (5'h7 == index_addr) begin // @[ICache.scala 110:26]
      if (update & updateway1) begin // @[ICache.scala 110:32]
        block1_7 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 64:39]
        block1_7 <= block1_31; // @[ICache.scala 64:39]
      end else begin
        block1_7 <= _GEN_159;
      end
    end
    if (reset) begin // @[ICache.scala 56:26]
      block1_8 <= 512'h0; // @[ICache.scala 56:26]
    end else if (5'h8 == index_addr) begin // @[ICache.scala 110:26]
      if (update & updateway1) begin // @[ICache.scala 110:32]
        block1_8 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 64:39]
        block1_8 <= block1_31; // @[ICache.scala 64:39]
      end else begin
        block1_8 <= _GEN_159;
      end
    end
    if (reset) begin // @[ICache.scala 56:26]
      block1_9 <= 512'h0; // @[ICache.scala 56:26]
    end else if (5'h9 == index_addr) begin // @[ICache.scala 110:26]
      if (update & updateway1) begin // @[ICache.scala 110:32]
        block1_9 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 64:39]
        block1_9 <= block1_31; // @[ICache.scala 64:39]
      end else begin
        block1_9 <= _GEN_159;
      end
    end
    if (reset) begin // @[ICache.scala 56:26]
      block1_10 <= 512'h0; // @[ICache.scala 56:26]
    end else if (5'ha == index_addr) begin // @[ICache.scala 110:26]
      if (update & updateway1) begin // @[ICache.scala 110:32]
        block1_10 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 64:39]
        block1_10 <= block1_31; // @[ICache.scala 64:39]
      end else begin
        block1_10 <= _GEN_159;
      end
    end
    if (reset) begin // @[ICache.scala 56:26]
      block1_11 <= 512'h0; // @[ICache.scala 56:26]
    end else if (5'hb == index_addr) begin // @[ICache.scala 110:26]
      if (update & updateway1) begin // @[ICache.scala 110:32]
        block1_11 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 64:39]
        block1_11 <= block1_31; // @[ICache.scala 64:39]
      end else begin
        block1_11 <= _GEN_159;
      end
    end
    if (reset) begin // @[ICache.scala 56:26]
      block1_12 <= 512'h0; // @[ICache.scala 56:26]
    end else if (5'hc == index_addr) begin // @[ICache.scala 110:26]
      if (update & updateway1) begin // @[ICache.scala 110:32]
        block1_12 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 64:39]
        block1_12 <= block1_31; // @[ICache.scala 64:39]
      end else begin
        block1_12 <= _GEN_159;
      end
    end
    if (reset) begin // @[ICache.scala 56:26]
      block1_13 <= 512'h0; // @[ICache.scala 56:26]
    end else if (5'hd == index_addr) begin // @[ICache.scala 110:26]
      if (update & updateway1) begin // @[ICache.scala 110:32]
        block1_13 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 64:39]
        block1_13 <= block1_31; // @[ICache.scala 64:39]
      end else begin
        block1_13 <= _GEN_159;
      end
    end
    if (reset) begin // @[ICache.scala 56:26]
      block1_14 <= 512'h0; // @[ICache.scala 56:26]
    end else if (5'he == index_addr) begin // @[ICache.scala 110:26]
      if (update & updateway1) begin // @[ICache.scala 110:32]
        block1_14 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 64:39]
        block1_14 <= block1_31; // @[ICache.scala 64:39]
      end else begin
        block1_14 <= _GEN_159;
      end
    end
    if (reset) begin // @[ICache.scala 56:26]
      block1_15 <= 512'h0; // @[ICache.scala 56:26]
    end else if (5'hf == index_addr) begin // @[ICache.scala 110:26]
      if (update & updateway1) begin // @[ICache.scala 110:32]
        block1_15 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 64:39]
        block1_15 <= block1_31; // @[ICache.scala 64:39]
      end else begin
        block1_15 <= _GEN_159;
      end
    end
    if (reset) begin // @[ICache.scala 56:26]
      block1_16 <= 512'h0; // @[ICache.scala 56:26]
    end else if (5'h10 == index_addr) begin // @[ICache.scala 110:26]
      if (update & updateway1) begin // @[ICache.scala 110:32]
        block1_16 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 64:39]
        block1_16 <= block1_31; // @[ICache.scala 64:39]
      end else begin
        block1_16 <= _GEN_159;
      end
    end
    if (reset) begin // @[ICache.scala 56:26]
      block1_17 <= 512'h0; // @[ICache.scala 56:26]
    end else if (5'h11 == index_addr) begin // @[ICache.scala 110:26]
      if (update & updateway1) begin // @[ICache.scala 110:32]
        block1_17 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 64:39]
        block1_17 <= block1_31; // @[ICache.scala 64:39]
      end else begin
        block1_17 <= _GEN_159;
      end
    end
    if (reset) begin // @[ICache.scala 56:26]
      block1_18 <= 512'h0; // @[ICache.scala 56:26]
    end else if (5'h12 == index_addr) begin // @[ICache.scala 110:26]
      if (update & updateway1) begin // @[ICache.scala 110:32]
        block1_18 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 64:39]
        block1_18 <= block1_31; // @[ICache.scala 64:39]
      end else begin
        block1_18 <= _GEN_159;
      end
    end
    if (reset) begin // @[ICache.scala 56:26]
      block1_19 <= 512'h0; // @[ICache.scala 56:26]
    end else if (5'h13 == index_addr) begin // @[ICache.scala 110:26]
      if (update & updateway1) begin // @[ICache.scala 110:32]
        block1_19 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 64:39]
        block1_19 <= block1_31; // @[ICache.scala 64:39]
      end else begin
        block1_19 <= _GEN_159;
      end
    end
    if (reset) begin // @[ICache.scala 56:26]
      block1_20 <= 512'h0; // @[ICache.scala 56:26]
    end else if (5'h14 == index_addr) begin // @[ICache.scala 110:26]
      if (update & updateway1) begin // @[ICache.scala 110:32]
        block1_20 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 64:39]
        block1_20 <= block1_31; // @[ICache.scala 64:39]
      end else begin
        block1_20 <= _GEN_159;
      end
    end
    if (reset) begin // @[ICache.scala 56:26]
      block1_21 <= 512'h0; // @[ICache.scala 56:26]
    end else if (5'h15 == index_addr) begin // @[ICache.scala 110:26]
      if (update & updateway1) begin // @[ICache.scala 110:32]
        block1_21 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 64:39]
        block1_21 <= block1_31; // @[ICache.scala 64:39]
      end else begin
        block1_21 <= _GEN_159;
      end
    end
    if (reset) begin // @[ICache.scala 56:26]
      block1_22 <= 512'h0; // @[ICache.scala 56:26]
    end else if (5'h16 == index_addr) begin // @[ICache.scala 110:26]
      if (update & updateway1) begin // @[ICache.scala 110:32]
        block1_22 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 64:39]
        block1_22 <= block1_31; // @[ICache.scala 64:39]
      end else begin
        block1_22 <= _GEN_159;
      end
    end
    if (reset) begin // @[ICache.scala 56:26]
      block1_23 <= 512'h0; // @[ICache.scala 56:26]
    end else if (5'h17 == index_addr) begin // @[ICache.scala 110:26]
      if (update & updateway1) begin // @[ICache.scala 110:32]
        block1_23 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 64:39]
        block1_23 <= block1_31; // @[ICache.scala 64:39]
      end else begin
        block1_23 <= _GEN_159;
      end
    end
    if (reset) begin // @[ICache.scala 56:26]
      block1_24 <= 512'h0; // @[ICache.scala 56:26]
    end else if (5'h18 == index_addr) begin // @[ICache.scala 110:26]
      if (update & updateway1) begin // @[ICache.scala 110:32]
        block1_24 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 64:39]
        block1_24 <= block1_31; // @[ICache.scala 64:39]
      end else begin
        block1_24 <= _GEN_159;
      end
    end
    if (reset) begin // @[ICache.scala 56:26]
      block1_25 <= 512'h0; // @[ICache.scala 56:26]
    end else if (5'h19 == index_addr) begin // @[ICache.scala 110:26]
      if (update & updateway1) begin // @[ICache.scala 110:32]
        block1_25 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 64:39]
        block1_25 <= block1_31; // @[ICache.scala 64:39]
      end else begin
        block1_25 <= _GEN_159;
      end
    end
    if (reset) begin // @[ICache.scala 56:26]
      block1_26 <= 512'h0; // @[ICache.scala 56:26]
    end else if (5'h1a == index_addr) begin // @[ICache.scala 110:26]
      if (update & updateway1) begin // @[ICache.scala 110:32]
        block1_26 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 64:39]
        block1_26 <= block1_31; // @[ICache.scala 64:39]
      end else begin
        block1_26 <= _GEN_159;
      end
    end
    if (reset) begin // @[ICache.scala 56:26]
      block1_27 <= 512'h0; // @[ICache.scala 56:26]
    end else if (5'h1b == index_addr) begin // @[ICache.scala 110:26]
      if (update & updateway1) begin // @[ICache.scala 110:32]
        block1_27 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 64:39]
        block1_27 <= block1_31; // @[ICache.scala 64:39]
      end else begin
        block1_27 <= _GEN_159;
      end
    end
    if (reset) begin // @[ICache.scala 56:26]
      block1_28 <= 512'h0; // @[ICache.scala 56:26]
    end else if (5'h1c == index_addr) begin // @[ICache.scala 110:26]
      if (update & updateway1) begin // @[ICache.scala 110:32]
        block1_28 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 64:39]
        block1_28 <= block1_31; // @[ICache.scala 64:39]
      end else begin
        block1_28 <= _GEN_159;
      end
    end
    if (reset) begin // @[ICache.scala 56:26]
      block1_29 <= 512'h0; // @[ICache.scala 56:26]
    end else if (5'h1d == index_addr) begin // @[ICache.scala 110:26]
      if (update & updateway1) begin // @[ICache.scala 110:32]
        block1_29 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 64:39]
        block1_29 <= block1_31; // @[ICache.scala 64:39]
      end else begin
        block1_29 <= _GEN_159;
      end
    end
    if (reset) begin // @[ICache.scala 56:26]
      block1_30 <= 512'h0; // @[ICache.scala 56:26]
    end else if (5'h1e == index_addr) begin // @[ICache.scala 110:26]
      if (update & updateway1) begin // @[ICache.scala 110:32]
        block1_30 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 64:39]
        block1_30 <= block1_31; // @[ICache.scala 64:39]
      end else begin
        block1_30 <= _GEN_159;
      end
    end
    if (reset) begin // @[ICache.scala 56:26]
      block1_31 <= 512'h0; // @[ICache.scala 56:26]
    end else if (5'h1f == index_addr) begin // @[ICache.scala 110:26]
      if (update & updateway1) begin // @[ICache.scala 110:32]
        block1_31 <= io_axi_data;
      end else if (!(5'h1f == index_addr)) begin // @[ICache.scala 64:39]
        block1_31 <= _GEN_159;
      end
    end
    if (reset) begin // @[ICache.scala 57:26]
      v2_0 <= 1'h0; // @[ICache.scala 57:26]
    end else if (state == 2'h3) begin // @[ICache.scala 119:37]
      if (5'h0 == fence_cnt) begin // @[ICache.scala 119:52]
        v2_0 <= 1'h0; // @[ICache.scala 119:52]
      end else begin
        v2_0 <= _GEN_490;
      end
    end else if (_block2_T) begin // @[ICache.scala 120:37]
      v2_0 <= _GEN_779 | _GEN_490;
    end else begin
      v2_0 <= _GEN_490;
    end
    if (reset) begin // @[ICache.scala 57:26]
      v2_1 <= 1'h0; // @[ICache.scala 57:26]
    end else if (state == 2'h3) begin // @[ICache.scala 119:37]
      if (5'h1 == fence_cnt) begin // @[ICache.scala 119:52]
        v2_1 <= 1'h0; // @[ICache.scala 119:52]
      end else begin
        v2_1 <= _GEN_491;
      end
    end else if (_block2_T) begin // @[ICache.scala 120:37]
      v2_1 <= _GEN_780 | _GEN_491;
    end else begin
      v2_1 <= _GEN_491;
    end
    if (reset) begin // @[ICache.scala 57:26]
      v2_2 <= 1'h0; // @[ICache.scala 57:26]
    end else if (state == 2'h3) begin // @[ICache.scala 119:37]
      if (5'h2 == fence_cnt) begin // @[ICache.scala 119:52]
        v2_2 <= 1'h0; // @[ICache.scala 119:52]
      end else begin
        v2_2 <= _GEN_492;
      end
    end else if (_block2_T) begin // @[ICache.scala 120:37]
      v2_2 <= _GEN_781 | _GEN_492;
    end else begin
      v2_2 <= _GEN_492;
    end
    if (reset) begin // @[ICache.scala 57:26]
      v2_3 <= 1'h0; // @[ICache.scala 57:26]
    end else if (state == 2'h3) begin // @[ICache.scala 119:37]
      if (5'h3 == fence_cnt) begin // @[ICache.scala 119:52]
        v2_3 <= 1'h0; // @[ICache.scala 119:52]
      end else begin
        v2_3 <= _GEN_493;
      end
    end else if (_block2_T) begin // @[ICache.scala 120:37]
      v2_3 <= _GEN_782 | _GEN_493;
    end else begin
      v2_3 <= _GEN_493;
    end
    if (reset) begin // @[ICache.scala 57:26]
      v2_4 <= 1'h0; // @[ICache.scala 57:26]
    end else if (state == 2'h3) begin // @[ICache.scala 119:37]
      if (5'h4 == fence_cnt) begin // @[ICache.scala 119:52]
        v2_4 <= 1'h0; // @[ICache.scala 119:52]
      end else begin
        v2_4 <= _GEN_494;
      end
    end else if (_block2_T) begin // @[ICache.scala 120:37]
      v2_4 <= _GEN_783 | _GEN_494;
    end else begin
      v2_4 <= _GEN_494;
    end
    if (reset) begin // @[ICache.scala 57:26]
      v2_5 <= 1'h0; // @[ICache.scala 57:26]
    end else if (state == 2'h3) begin // @[ICache.scala 119:37]
      if (5'h5 == fence_cnt) begin // @[ICache.scala 119:52]
        v2_5 <= 1'h0; // @[ICache.scala 119:52]
      end else begin
        v2_5 <= _GEN_495;
      end
    end else if (_block2_T) begin // @[ICache.scala 120:37]
      v2_5 <= _GEN_784 | _GEN_495;
    end else begin
      v2_5 <= _GEN_495;
    end
    if (reset) begin // @[ICache.scala 57:26]
      v2_6 <= 1'h0; // @[ICache.scala 57:26]
    end else if (state == 2'h3) begin // @[ICache.scala 119:37]
      if (5'h6 == fence_cnt) begin // @[ICache.scala 119:52]
        v2_6 <= 1'h0; // @[ICache.scala 119:52]
      end else begin
        v2_6 <= _GEN_496;
      end
    end else if (_block2_T) begin // @[ICache.scala 120:37]
      v2_6 <= _GEN_785 | _GEN_496;
    end else begin
      v2_6 <= _GEN_496;
    end
    if (reset) begin // @[ICache.scala 57:26]
      v2_7 <= 1'h0; // @[ICache.scala 57:26]
    end else if (state == 2'h3) begin // @[ICache.scala 119:37]
      if (5'h7 == fence_cnt) begin // @[ICache.scala 119:52]
        v2_7 <= 1'h0; // @[ICache.scala 119:52]
      end else begin
        v2_7 <= _GEN_497;
      end
    end else if (_block2_T) begin // @[ICache.scala 120:37]
      v2_7 <= _GEN_786 | _GEN_497;
    end else begin
      v2_7 <= _GEN_497;
    end
    if (reset) begin // @[ICache.scala 57:26]
      v2_8 <= 1'h0; // @[ICache.scala 57:26]
    end else if (state == 2'h3) begin // @[ICache.scala 119:37]
      if (5'h8 == fence_cnt) begin // @[ICache.scala 119:52]
        v2_8 <= 1'h0; // @[ICache.scala 119:52]
      end else begin
        v2_8 <= _GEN_498;
      end
    end else if (_block2_T) begin // @[ICache.scala 120:37]
      v2_8 <= _GEN_787 | _GEN_498;
    end else begin
      v2_8 <= _GEN_498;
    end
    if (reset) begin // @[ICache.scala 57:26]
      v2_9 <= 1'h0; // @[ICache.scala 57:26]
    end else if (state == 2'h3) begin // @[ICache.scala 119:37]
      if (5'h9 == fence_cnt) begin // @[ICache.scala 119:52]
        v2_9 <= 1'h0; // @[ICache.scala 119:52]
      end else begin
        v2_9 <= _GEN_499;
      end
    end else if (_block2_T) begin // @[ICache.scala 120:37]
      v2_9 <= _GEN_788 | _GEN_499;
    end else begin
      v2_9 <= _GEN_499;
    end
    if (reset) begin // @[ICache.scala 57:26]
      v2_10 <= 1'h0; // @[ICache.scala 57:26]
    end else if (state == 2'h3) begin // @[ICache.scala 119:37]
      if (5'ha == fence_cnt) begin // @[ICache.scala 119:52]
        v2_10 <= 1'h0; // @[ICache.scala 119:52]
      end else begin
        v2_10 <= _GEN_500;
      end
    end else if (_block2_T) begin // @[ICache.scala 120:37]
      v2_10 <= _GEN_789 | _GEN_500;
    end else begin
      v2_10 <= _GEN_500;
    end
    if (reset) begin // @[ICache.scala 57:26]
      v2_11 <= 1'h0; // @[ICache.scala 57:26]
    end else if (state == 2'h3) begin // @[ICache.scala 119:37]
      if (5'hb == fence_cnt) begin // @[ICache.scala 119:52]
        v2_11 <= 1'h0; // @[ICache.scala 119:52]
      end else begin
        v2_11 <= _GEN_501;
      end
    end else if (_block2_T) begin // @[ICache.scala 120:37]
      v2_11 <= _GEN_790 | _GEN_501;
    end else begin
      v2_11 <= _GEN_501;
    end
    if (reset) begin // @[ICache.scala 57:26]
      v2_12 <= 1'h0; // @[ICache.scala 57:26]
    end else if (state == 2'h3) begin // @[ICache.scala 119:37]
      if (5'hc == fence_cnt) begin // @[ICache.scala 119:52]
        v2_12 <= 1'h0; // @[ICache.scala 119:52]
      end else begin
        v2_12 <= _GEN_502;
      end
    end else if (_block2_T) begin // @[ICache.scala 120:37]
      v2_12 <= _GEN_791 | _GEN_502;
    end else begin
      v2_12 <= _GEN_502;
    end
    if (reset) begin // @[ICache.scala 57:26]
      v2_13 <= 1'h0; // @[ICache.scala 57:26]
    end else if (state == 2'h3) begin // @[ICache.scala 119:37]
      if (5'hd == fence_cnt) begin // @[ICache.scala 119:52]
        v2_13 <= 1'h0; // @[ICache.scala 119:52]
      end else begin
        v2_13 <= _GEN_503;
      end
    end else if (_block2_T) begin // @[ICache.scala 120:37]
      v2_13 <= _GEN_792 | _GEN_503;
    end else begin
      v2_13 <= _GEN_503;
    end
    if (reset) begin // @[ICache.scala 57:26]
      v2_14 <= 1'h0; // @[ICache.scala 57:26]
    end else if (state == 2'h3) begin // @[ICache.scala 119:37]
      if (5'he == fence_cnt) begin // @[ICache.scala 119:52]
        v2_14 <= 1'h0; // @[ICache.scala 119:52]
      end else begin
        v2_14 <= _GEN_504;
      end
    end else if (_block2_T) begin // @[ICache.scala 120:37]
      v2_14 <= _GEN_793 | _GEN_504;
    end else begin
      v2_14 <= _GEN_504;
    end
    if (reset) begin // @[ICache.scala 57:26]
      v2_15 <= 1'h0; // @[ICache.scala 57:26]
    end else if (state == 2'h3) begin // @[ICache.scala 119:37]
      if (5'hf == fence_cnt) begin // @[ICache.scala 119:52]
        v2_15 <= 1'h0; // @[ICache.scala 119:52]
      end else begin
        v2_15 <= _GEN_505;
      end
    end else if (_block2_T) begin // @[ICache.scala 120:37]
      v2_15 <= _GEN_794 | _GEN_505;
    end else begin
      v2_15 <= _GEN_505;
    end
    if (reset) begin // @[ICache.scala 57:26]
      v2_16 <= 1'h0; // @[ICache.scala 57:26]
    end else if (state == 2'h3) begin // @[ICache.scala 119:37]
      if (5'h10 == fence_cnt) begin // @[ICache.scala 119:52]
        v2_16 <= 1'h0; // @[ICache.scala 119:52]
      end else begin
        v2_16 <= _GEN_506;
      end
    end else if (_block2_T) begin // @[ICache.scala 120:37]
      v2_16 <= _GEN_795 | _GEN_506;
    end else begin
      v2_16 <= _GEN_506;
    end
    if (reset) begin // @[ICache.scala 57:26]
      v2_17 <= 1'h0; // @[ICache.scala 57:26]
    end else if (state == 2'h3) begin // @[ICache.scala 119:37]
      if (5'h11 == fence_cnt) begin // @[ICache.scala 119:52]
        v2_17 <= 1'h0; // @[ICache.scala 119:52]
      end else begin
        v2_17 <= _GEN_507;
      end
    end else if (_block2_T) begin // @[ICache.scala 120:37]
      v2_17 <= _GEN_796 | _GEN_507;
    end else begin
      v2_17 <= _GEN_507;
    end
    if (reset) begin // @[ICache.scala 57:26]
      v2_18 <= 1'h0; // @[ICache.scala 57:26]
    end else if (state == 2'h3) begin // @[ICache.scala 119:37]
      if (5'h12 == fence_cnt) begin // @[ICache.scala 119:52]
        v2_18 <= 1'h0; // @[ICache.scala 119:52]
      end else begin
        v2_18 <= _GEN_508;
      end
    end else if (_block2_T) begin // @[ICache.scala 120:37]
      v2_18 <= _GEN_797 | _GEN_508;
    end else begin
      v2_18 <= _GEN_508;
    end
    if (reset) begin // @[ICache.scala 57:26]
      v2_19 <= 1'h0; // @[ICache.scala 57:26]
    end else if (state == 2'h3) begin // @[ICache.scala 119:37]
      if (5'h13 == fence_cnt) begin // @[ICache.scala 119:52]
        v2_19 <= 1'h0; // @[ICache.scala 119:52]
      end else begin
        v2_19 <= _GEN_509;
      end
    end else if (_block2_T) begin // @[ICache.scala 120:37]
      v2_19 <= _GEN_798 | _GEN_509;
    end else begin
      v2_19 <= _GEN_509;
    end
    if (reset) begin // @[ICache.scala 57:26]
      v2_20 <= 1'h0; // @[ICache.scala 57:26]
    end else if (state == 2'h3) begin // @[ICache.scala 119:37]
      if (5'h14 == fence_cnt) begin // @[ICache.scala 119:52]
        v2_20 <= 1'h0; // @[ICache.scala 119:52]
      end else begin
        v2_20 <= _GEN_510;
      end
    end else if (_block2_T) begin // @[ICache.scala 120:37]
      v2_20 <= _GEN_799 | _GEN_510;
    end else begin
      v2_20 <= _GEN_510;
    end
    if (reset) begin // @[ICache.scala 57:26]
      v2_21 <= 1'h0; // @[ICache.scala 57:26]
    end else if (state == 2'h3) begin // @[ICache.scala 119:37]
      if (5'h15 == fence_cnt) begin // @[ICache.scala 119:52]
        v2_21 <= 1'h0; // @[ICache.scala 119:52]
      end else begin
        v2_21 <= _GEN_511;
      end
    end else if (_block2_T) begin // @[ICache.scala 120:37]
      v2_21 <= _GEN_800 | _GEN_511;
    end else begin
      v2_21 <= _GEN_511;
    end
    if (reset) begin // @[ICache.scala 57:26]
      v2_22 <= 1'h0; // @[ICache.scala 57:26]
    end else if (state == 2'h3) begin // @[ICache.scala 119:37]
      if (5'h16 == fence_cnt) begin // @[ICache.scala 119:52]
        v2_22 <= 1'h0; // @[ICache.scala 119:52]
      end else begin
        v2_22 <= _GEN_512;
      end
    end else if (_block2_T) begin // @[ICache.scala 120:37]
      v2_22 <= _GEN_801 | _GEN_512;
    end else begin
      v2_22 <= _GEN_512;
    end
    if (reset) begin // @[ICache.scala 57:26]
      v2_23 <= 1'h0; // @[ICache.scala 57:26]
    end else if (state == 2'h3) begin // @[ICache.scala 119:37]
      if (5'h17 == fence_cnt) begin // @[ICache.scala 119:52]
        v2_23 <= 1'h0; // @[ICache.scala 119:52]
      end else begin
        v2_23 <= _GEN_513;
      end
    end else if (_block2_T) begin // @[ICache.scala 120:37]
      v2_23 <= _GEN_802 | _GEN_513;
    end else begin
      v2_23 <= _GEN_513;
    end
    if (reset) begin // @[ICache.scala 57:26]
      v2_24 <= 1'h0; // @[ICache.scala 57:26]
    end else if (state == 2'h3) begin // @[ICache.scala 119:37]
      if (5'h18 == fence_cnt) begin // @[ICache.scala 119:52]
        v2_24 <= 1'h0; // @[ICache.scala 119:52]
      end else begin
        v2_24 <= _GEN_514;
      end
    end else if (_block2_T) begin // @[ICache.scala 120:37]
      v2_24 <= _GEN_803 | _GEN_514;
    end else begin
      v2_24 <= _GEN_514;
    end
    if (reset) begin // @[ICache.scala 57:26]
      v2_25 <= 1'h0; // @[ICache.scala 57:26]
    end else if (state == 2'h3) begin // @[ICache.scala 119:37]
      if (5'h19 == fence_cnt) begin // @[ICache.scala 119:52]
        v2_25 <= 1'h0; // @[ICache.scala 119:52]
      end else begin
        v2_25 <= _GEN_515;
      end
    end else if (_block2_T) begin // @[ICache.scala 120:37]
      v2_25 <= _GEN_804 | _GEN_515;
    end else begin
      v2_25 <= _GEN_515;
    end
    if (reset) begin // @[ICache.scala 57:26]
      v2_26 <= 1'h0; // @[ICache.scala 57:26]
    end else if (state == 2'h3) begin // @[ICache.scala 119:37]
      if (5'h1a == fence_cnt) begin // @[ICache.scala 119:52]
        v2_26 <= 1'h0; // @[ICache.scala 119:52]
      end else begin
        v2_26 <= _GEN_516;
      end
    end else if (_block2_T) begin // @[ICache.scala 120:37]
      v2_26 <= _GEN_805 | _GEN_516;
    end else begin
      v2_26 <= _GEN_516;
    end
    if (reset) begin // @[ICache.scala 57:26]
      v2_27 <= 1'h0; // @[ICache.scala 57:26]
    end else if (state == 2'h3) begin // @[ICache.scala 119:37]
      if (5'h1b == fence_cnt) begin // @[ICache.scala 119:52]
        v2_27 <= 1'h0; // @[ICache.scala 119:52]
      end else begin
        v2_27 <= _GEN_517;
      end
    end else if (_block2_T) begin // @[ICache.scala 120:37]
      v2_27 <= _GEN_806 | _GEN_517;
    end else begin
      v2_27 <= _GEN_517;
    end
    if (reset) begin // @[ICache.scala 57:26]
      v2_28 <= 1'h0; // @[ICache.scala 57:26]
    end else if (state == 2'h3) begin // @[ICache.scala 119:37]
      if (5'h1c == fence_cnt) begin // @[ICache.scala 119:52]
        v2_28 <= 1'h0; // @[ICache.scala 119:52]
      end else begin
        v2_28 <= _GEN_518;
      end
    end else if (_block2_T) begin // @[ICache.scala 120:37]
      v2_28 <= _GEN_807 | _GEN_518;
    end else begin
      v2_28 <= _GEN_518;
    end
    if (reset) begin // @[ICache.scala 57:26]
      v2_29 <= 1'h0; // @[ICache.scala 57:26]
    end else if (state == 2'h3) begin // @[ICache.scala 119:37]
      if (5'h1d == fence_cnt) begin // @[ICache.scala 119:52]
        v2_29 <= 1'h0; // @[ICache.scala 119:52]
      end else begin
        v2_29 <= _GEN_519;
      end
    end else if (_block2_T) begin // @[ICache.scala 120:37]
      v2_29 <= _GEN_808 | _GEN_519;
    end else begin
      v2_29 <= _GEN_519;
    end
    if (reset) begin // @[ICache.scala 57:26]
      v2_30 <= 1'h0; // @[ICache.scala 57:26]
    end else if (state == 2'h3) begin // @[ICache.scala 119:37]
      if (5'h1e == fence_cnt) begin // @[ICache.scala 119:52]
        v2_30 <= 1'h0; // @[ICache.scala 119:52]
      end else begin
        v2_30 <= _GEN_520;
      end
    end else if (_block2_T) begin // @[ICache.scala 120:37]
      v2_30 <= _GEN_809 | _GEN_520;
    end else begin
      v2_30 <= _GEN_520;
    end
    if (reset) begin // @[ICache.scala 57:26]
      v2_31 <= 1'h0; // @[ICache.scala 57:26]
    end else if (state == 2'h3) begin // @[ICache.scala 119:37]
      if (5'h1f == fence_cnt) begin // @[ICache.scala 119:52]
        v2_31 <= 1'h0; // @[ICache.scala 119:52]
      end else begin
        v2_31 <= _GEN_521;
      end
    end else if (_block2_T) begin // @[ICache.scala 120:37]
      v2_31 <= _GEN_810 | _GEN_521;
    end else begin
      v2_31 <= _GEN_521;
    end
    if (reset) begin // @[ICache.scala 58:26]
      age2_0 <= 1'h0; // @[ICache.scala 58:26]
    end else if (5'h0 == index_addr) begin // @[ICache.scala 72:22]
      if (_age1_T) begin // @[ICache.scala 72:28]
        age2_0 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 72:28]
        age2_0 <= age2_31; // @[ICache.scala 72:28]
      end else begin
        age2_0 <= _GEN_287;
      end
    end
    if (reset) begin // @[ICache.scala 58:26]
      age2_1 <= 1'h0; // @[ICache.scala 58:26]
    end else if (5'h1 == index_addr) begin // @[ICache.scala 72:22]
      if (_age1_T) begin // @[ICache.scala 72:28]
        age2_1 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 72:28]
        age2_1 <= age2_31; // @[ICache.scala 72:28]
      end else begin
        age2_1 <= _GEN_287;
      end
    end
    if (reset) begin // @[ICache.scala 58:26]
      age2_2 <= 1'h0; // @[ICache.scala 58:26]
    end else if (5'h2 == index_addr) begin // @[ICache.scala 72:22]
      if (_age1_T) begin // @[ICache.scala 72:28]
        age2_2 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 72:28]
        age2_2 <= age2_31; // @[ICache.scala 72:28]
      end else begin
        age2_2 <= _GEN_287;
      end
    end
    if (reset) begin // @[ICache.scala 58:26]
      age2_3 <= 1'h0; // @[ICache.scala 58:26]
    end else if (5'h3 == index_addr) begin // @[ICache.scala 72:22]
      if (_age1_T) begin // @[ICache.scala 72:28]
        age2_3 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 72:28]
        age2_3 <= age2_31; // @[ICache.scala 72:28]
      end else begin
        age2_3 <= _GEN_287;
      end
    end
    if (reset) begin // @[ICache.scala 58:26]
      age2_4 <= 1'h0; // @[ICache.scala 58:26]
    end else if (5'h4 == index_addr) begin // @[ICache.scala 72:22]
      if (_age1_T) begin // @[ICache.scala 72:28]
        age2_4 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 72:28]
        age2_4 <= age2_31; // @[ICache.scala 72:28]
      end else begin
        age2_4 <= _GEN_287;
      end
    end
    if (reset) begin // @[ICache.scala 58:26]
      age2_5 <= 1'h0; // @[ICache.scala 58:26]
    end else if (5'h5 == index_addr) begin // @[ICache.scala 72:22]
      if (_age1_T) begin // @[ICache.scala 72:28]
        age2_5 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 72:28]
        age2_5 <= age2_31; // @[ICache.scala 72:28]
      end else begin
        age2_5 <= _GEN_287;
      end
    end
    if (reset) begin // @[ICache.scala 58:26]
      age2_6 <= 1'h0; // @[ICache.scala 58:26]
    end else if (5'h6 == index_addr) begin // @[ICache.scala 72:22]
      if (_age1_T) begin // @[ICache.scala 72:28]
        age2_6 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 72:28]
        age2_6 <= age2_31; // @[ICache.scala 72:28]
      end else begin
        age2_6 <= _GEN_287;
      end
    end
    if (reset) begin // @[ICache.scala 58:26]
      age2_7 <= 1'h0; // @[ICache.scala 58:26]
    end else if (5'h7 == index_addr) begin // @[ICache.scala 72:22]
      if (_age1_T) begin // @[ICache.scala 72:28]
        age2_7 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 72:28]
        age2_7 <= age2_31; // @[ICache.scala 72:28]
      end else begin
        age2_7 <= _GEN_287;
      end
    end
    if (reset) begin // @[ICache.scala 58:26]
      age2_8 <= 1'h0; // @[ICache.scala 58:26]
    end else if (5'h8 == index_addr) begin // @[ICache.scala 72:22]
      if (_age1_T) begin // @[ICache.scala 72:28]
        age2_8 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 72:28]
        age2_8 <= age2_31; // @[ICache.scala 72:28]
      end else begin
        age2_8 <= _GEN_287;
      end
    end
    if (reset) begin // @[ICache.scala 58:26]
      age2_9 <= 1'h0; // @[ICache.scala 58:26]
    end else if (5'h9 == index_addr) begin // @[ICache.scala 72:22]
      if (_age1_T) begin // @[ICache.scala 72:28]
        age2_9 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 72:28]
        age2_9 <= age2_31; // @[ICache.scala 72:28]
      end else begin
        age2_9 <= _GEN_287;
      end
    end
    if (reset) begin // @[ICache.scala 58:26]
      age2_10 <= 1'h0; // @[ICache.scala 58:26]
    end else if (5'ha == index_addr) begin // @[ICache.scala 72:22]
      if (_age1_T) begin // @[ICache.scala 72:28]
        age2_10 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 72:28]
        age2_10 <= age2_31; // @[ICache.scala 72:28]
      end else begin
        age2_10 <= _GEN_287;
      end
    end
    if (reset) begin // @[ICache.scala 58:26]
      age2_11 <= 1'h0; // @[ICache.scala 58:26]
    end else if (5'hb == index_addr) begin // @[ICache.scala 72:22]
      if (_age1_T) begin // @[ICache.scala 72:28]
        age2_11 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 72:28]
        age2_11 <= age2_31; // @[ICache.scala 72:28]
      end else begin
        age2_11 <= _GEN_287;
      end
    end
    if (reset) begin // @[ICache.scala 58:26]
      age2_12 <= 1'h0; // @[ICache.scala 58:26]
    end else if (5'hc == index_addr) begin // @[ICache.scala 72:22]
      if (_age1_T) begin // @[ICache.scala 72:28]
        age2_12 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 72:28]
        age2_12 <= age2_31; // @[ICache.scala 72:28]
      end else begin
        age2_12 <= _GEN_287;
      end
    end
    if (reset) begin // @[ICache.scala 58:26]
      age2_13 <= 1'h0; // @[ICache.scala 58:26]
    end else if (5'hd == index_addr) begin // @[ICache.scala 72:22]
      if (_age1_T) begin // @[ICache.scala 72:28]
        age2_13 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 72:28]
        age2_13 <= age2_31; // @[ICache.scala 72:28]
      end else begin
        age2_13 <= _GEN_287;
      end
    end
    if (reset) begin // @[ICache.scala 58:26]
      age2_14 <= 1'h0; // @[ICache.scala 58:26]
    end else if (5'he == index_addr) begin // @[ICache.scala 72:22]
      if (_age1_T) begin // @[ICache.scala 72:28]
        age2_14 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 72:28]
        age2_14 <= age2_31; // @[ICache.scala 72:28]
      end else begin
        age2_14 <= _GEN_287;
      end
    end
    if (reset) begin // @[ICache.scala 58:26]
      age2_15 <= 1'h0; // @[ICache.scala 58:26]
    end else if (5'hf == index_addr) begin // @[ICache.scala 72:22]
      if (_age1_T) begin // @[ICache.scala 72:28]
        age2_15 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 72:28]
        age2_15 <= age2_31; // @[ICache.scala 72:28]
      end else begin
        age2_15 <= _GEN_287;
      end
    end
    if (reset) begin // @[ICache.scala 58:26]
      age2_16 <= 1'h0; // @[ICache.scala 58:26]
    end else if (5'h10 == index_addr) begin // @[ICache.scala 72:22]
      if (_age1_T) begin // @[ICache.scala 72:28]
        age2_16 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 72:28]
        age2_16 <= age2_31; // @[ICache.scala 72:28]
      end else begin
        age2_16 <= _GEN_287;
      end
    end
    if (reset) begin // @[ICache.scala 58:26]
      age2_17 <= 1'h0; // @[ICache.scala 58:26]
    end else if (5'h11 == index_addr) begin // @[ICache.scala 72:22]
      if (_age1_T) begin // @[ICache.scala 72:28]
        age2_17 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 72:28]
        age2_17 <= age2_31; // @[ICache.scala 72:28]
      end else begin
        age2_17 <= _GEN_287;
      end
    end
    if (reset) begin // @[ICache.scala 58:26]
      age2_18 <= 1'h0; // @[ICache.scala 58:26]
    end else if (5'h12 == index_addr) begin // @[ICache.scala 72:22]
      if (_age1_T) begin // @[ICache.scala 72:28]
        age2_18 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 72:28]
        age2_18 <= age2_31; // @[ICache.scala 72:28]
      end else begin
        age2_18 <= _GEN_287;
      end
    end
    if (reset) begin // @[ICache.scala 58:26]
      age2_19 <= 1'h0; // @[ICache.scala 58:26]
    end else if (5'h13 == index_addr) begin // @[ICache.scala 72:22]
      if (_age1_T) begin // @[ICache.scala 72:28]
        age2_19 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 72:28]
        age2_19 <= age2_31; // @[ICache.scala 72:28]
      end else begin
        age2_19 <= _GEN_287;
      end
    end
    if (reset) begin // @[ICache.scala 58:26]
      age2_20 <= 1'h0; // @[ICache.scala 58:26]
    end else if (5'h14 == index_addr) begin // @[ICache.scala 72:22]
      if (_age1_T) begin // @[ICache.scala 72:28]
        age2_20 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 72:28]
        age2_20 <= age2_31; // @[ICache.scala 72:28]
      end else begin
        age2_20 <= _GEN_287;
      end
    end
    if (reset) begin // @[ICache.scala 58:26]
      age2_21 <= 1'h0; // @[ICache.scala 58:26]
    end else if (5'h15 == index_addr) begin // @[ICache.scala 72:22]
      if (_age1_T) begin // @[ICache.scala 72:28]
        age2_21 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 72:28]
        age2_21 <= age2_31; // @[ICache.scala 72:28]
      end else begin
        age2_21 <= _GEN_287;
      end
    end
    if (reset) begin // @[ICache.scala 58:26]
      age2_22 <= 1'h0; // @[ICache.scala 58:26]
    end else if (5'h16 == index_addr) begin // @[ICache.scala 72:22]
      if (_age1_T) begin // @[ICache.scala 72:28]
        age2_22 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 72:28]
        age2_22 <= age2_31; // @[ICache.scala 72:28]
      end else begin
        age2_22 <= _GEN_287;
      end
    end
    if (reset) begin // @[ICache.scala 58:26]
      age2_23 <= 1'h0; // @[ICache.scala 58:26]
    end else if (5'h17 == index_addr) begin // @[ICache.scala 72:22]
      if (_age1_T) begin // @[ICache.scala 72:28]
        age2_23 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 72:28]
        age2_23 <= age2_31; // @[ICache.scala 72:28]
      end else begin
        age2_23 <= _GEN_287;
      end
    end
    if (reset) begin // @[ICache.scala 58:26]
      age2_24 <= 1'h0; // @[ICache.scala 58:26]
    end else if (5'h18 == index_addr) begin // @[ICache.scala 72:22]
      if (_age1_T) begin // @[ICache.scala 72:28]
        age2_24 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 72:28]
        age2_24 <= age2_31; // @[ICache.scala 72:28]
      end else begin
        age2_24 <= _GEN_287;
      end
    end
    if (reset) begin // @[ICache.scala 58:26]
      age2_25 <= 1'h0; // @[ICache.scala 58:26]
    end else if (5'h19 == index_addr) begin // @[ICache.scala 72:22]
      if (_age1_T) begin // @[ICache.scala 72:28]
        age2_25 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 72:28]
        age2_25 <= age2_31; // @[ICache.scala 72:28]
      end else begin
        age2_25 <= _GEN_287;
      end
    end
    if (reset) begin // @[ICache.scala 58:26]
      age2_26 <= 1'h0; // @[ICache.scala 58:26]
    end else if (5'h1a == index_addr) begin // @[ICache.scala 72:22]
      if (_age1_T) begin // @[ICache.scala 72:28]
        age2_26 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 72:28]
        age2_26 <= age2_31; // @[ICache.scala 72:28]
      end else begin
        age2_26 <= _GEN_287;
      end
    end
    if (reset) begin // @[ICache.scala 58:26]
      age2_27 <= 1'h0; // @[ICache.scala 58:26]
    end else if (5'h1b == index_addr) begin // @[ICache.scala 72:22]
      if (_age1_T) begin // @[ICache.scala 72:28]
        age2_27 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 72:28]
        age2_27 <= age2_31; // @[ICache.scala 72:28]
      end else begin
        age2_27 <= _GEN_287;
      end
    end
    if (reset) begin // @[ICache.scala 58:26]
      age2_28 <= 1'h0; // @[ICache.scala 58:26]
    end else if (5'h1c == index_addr) begin // @[ICache.scala 72:22]
      if (_age1_T) begin // @[ICache.scala 72:28]
        age2_28 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 72:28]
        age2_28 <= age2_31; // @[ICache.scala 72:28]
      end else begin
        age2_28 <= _GEN_287;
      end
    end
    if (reset) begin // @[ICache.scala 58:26]
      age2_29 <= 1'h0; // @[ICache.scala 58:26]
    end else if (5'h1d == index_addr) begin // @[ICache.scala 72:22]
      if (_age1_T) begin // @[ICache.scala 72:28]
        age2_29 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 72:28]
        age2_29 <= age2_31; // @[ICache.scala 72:28]
      end else begin
        age2_29 <= _GEN_287;
      end
    end
    if (reset) begin // @[ICache.scala 58:26]
      age2_30 <= 1'h0; // @[ICache.scala 58:26]
    end else if (5'h1e == index_addr) begin // @[ICache.scala 72:22]
      if (_age1_T) begin // @[ICache.scala 72:28]
        age2_30 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 72:28]
        age2_30 <= age2_31; // @[ICache.scala 72:28]
      end else begin
        age2_30 <= _GEN_287;
      end
    end
    if (reset) begin // @[ICache.scala 58:26]
      age2_31 <= 1'h0; // @[ICache.scala 58:26]
    end else if (5'h1f == index_addr) begin // @[ICache.scala 72:22]
      if (_age1_T) begin // @[ICache.scala 72:28]
        age2_31 <= hit2;
      end else if (!(5'h1f == index_addr)) begin // @[ICache.scala 72:28]
        age2_31 <= _GEN_287;
      end
    end
    if (reset) begin // @[ICache.scala 59:26]
      tag2_0 <= 53'h0; // @[ICache.scala 59:26]
    end else if (5'h0 == index_addr) begin // @[ICache.scala 114:26]
      if (_block2_T) begin // @[ICache.scala 114:32]
        tag2_0 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 63:28]
        tag2_0 <= tag2_31; // @[ICache.scala 63:28]
      end else begin
        tag2_0 <= _GEN_95;
      end
    end
    if (reset) begin // @[ICache.scala 59:26]
      tag2_1 <= 53'h0; // @[ICache.scala 59:26]
    end else if (5'h1 == index_addr) begin // @[ICache.scala 114:26]
      if (_block2_T) begin // @[ICache.scala 114:32]
        tag2_1 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 63:28]
        tag2_1 <= tag2_31; // @[ICache.scala 63:28]
      end else begin
        tag2_1 <= _GEN_95;
      end
    end
    if (reset) begin // @[ICache.scala 59:26]
      tag2_2 <= 53'h0; // @[ICache.scala 59:26]
    end else if (5'h2 == index_addr) begin // @[ICache.scala 114:26]
      if (_block2_T) begin // @[ICache.scala 114:32]
        tag2_2 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 63:28]
        tag2_2 <= tag2_31; // @[ICache.scala 63:28]
      end else begin
        tag2_2 <= _GEN_95;
      end
    end
    if (reset) begin // @[ICache.scala 59:26]
      tag2_3 <= 53'h0; // @[ICache.scala 59:26]
    end else if (5'h3 == index_addr) begin // @[ICache.scala 114:26]
      if (_block2_T) begin // @[ICache.scala 114:32]
        tag2_3 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 63:28]
        tag2_3 <= tag2_31; // @[ICache.scala 63:28]
      end else begin
        tag2_3 <= _GEN_95;
      end
    end
    if (reset) begin // @[ICache.scala 59:26]
      tag2_4 <= 53'h0; // @[ICache.scala 59:26]
    end else if (5'h4 == index_addr) begin // @[ICache.scala 114:26]
      if (_block2_T) begin // @[ICache.scala 114:32]
        tag2_4 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 63:28]
        tag2_4 <= tag2_31; // @[ICache.scala 63:28]
      end else begin
        tag2_4 <= _GEN_95;
      end
    end
    if (reset) begin // @[ICache.scala 59:26]
      tag2_5 <= 53'h0; // @[ICache.scala 59:26]
    end else if (5'h5 == index_addr) begin // @[ICache.scala 114:26]
      if (_block2_T) begin // @[ICache.scala 114:32]
        tag2_5 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 63:28]
        tag2_5 <= tag2_31; // @[ICache.scala 63:28]
      end else begin
        tag2_5 <= _GEN_95;
      end
    end
    if (reset) begin // @[ICache.scala 59:26]
      tag2_6 <= 53'h0; // @[ICache.scala 59:26]
    end else if (5'h6 == index_addr) begin // @[ICache.scala 114:26]
      if (_block2_T) begin // @[ICache.scala 114:32]
        tag2_6 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 63:28]
        tag2_6 <= tag2_31; // @[ICache.scala 63:28]
      end else begin
        tag2_6 <= _GEN_95;
      end
    end
    if (reset) begin // @[ICache.scala 59:26]
      tag2_7 <= 53'h0; // @[ICache.scala 59:26]
    end else if (5'h7 == index_addr) begin // @[ICache.scala 114:26]
      if (_block2_T) begin // @[ICache.scala 114:32]
        tag2_7 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 63:28]
        tag2_7 <= tag2_31; // @[ICache.scala 63:28]
      end else begin
        tag2_7 <= _GEN_95;
      end
    end
    if (reset) begin // @[ICache.scala 59:26]
      tag2_8 <= 53'h0; // @[ICache.scala 59:26]
    end else if (5'h8 == index_addr) begin // @[ICache.scala 114:26]
      if (_block2_T) begin // @[ICache.scala 114:32]
        tag2_8 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 63:28]
        tag2_8 <= tag2_31; // @[ICache.scala 63:28]
      end else begin
        tag2_8 <= _GEN_95;
      end
    end
    if (reset) begin // @[ICache.scala 59:26]
      tag2_9 <= 53'h0; // @[ICache.scala 59:26]
    end else if (5'h9 == index_addr) begin // @[ICache.scala 114:26]
      if (_block2_T) begin // @[ICache.scala 114:32]
        tag2_9 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 63:28]
        tag2_9 <= tag2_31; // @[ICache.scala 63:28]
      end else begin
        tag2_9 <= _GEN_95;
      end
    end
    if (reset) begin // @[ICache.scala 59:26]
      tag2_10 <= 53'h0; // @[ICache.scala 59:26]
    end else if (5'ha == index_addr) begin // @[ICache.scala 114:26]
      if (_block2_T) begin // @[ICache.scala 114:32]
        tag2_10 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 63:28]
        tag2_10 <= tag2_31; // @[ICache.scala 63:28]
      end else begin
        tag2_10 <= _GEN_95;
      end
    end
    if (reset) begin // @[ICache.scala 59:26]
      tag2_11 <= 53'h0; // @[ICache.scala 59:26]
    end else if (5'hb == index_addr) begin // @[ICache.scala 114:26]
      if (_block2_T) begin // @[ICache.scala 114:32]
        tag2_11 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 63:28]
        tag2_11 <= tag2_31; // @[ICache.scala 63:28]
      end else begin
        tag2_11 <= _GEN_95;
      end
    end
    if (reset) begin // @[ICache.scala 59:26]
      tag2_12 <= 53'h0; // @[ICache.scala 59:26]
    end else if (5'hc == index_addr) begin // @[ICache.scala 114:26]
      if (_block2_T) begin // @[ICache.scala 114:32]
        tag2_12 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 63:28]
        tag2_12 <= tag2_31; // @[ICache.scala 63:28]
      end else begin
        tag2_12 <= _GEN_95;
      end
    end
    if (reset) begin // @[ICache.scala 59:26]
      tag2_13 <= 53'h0; // @[ICache.scala 59:26]
    end else if (5'hd == index_addr) begin // @[ICache.scala 114:26]
      if (_block2_T) begin // @[ICache.scala 114:32]
        tag2_13 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 63:28]
        tag2_13 <= tag2_31; // @[ICache.scala 63:28]
      end else begin
        tag2_13 <= _GEN_95;
      end
    end
    if (reset) begin // @[ICache.scala 59:26]
      tag2_14 <= 53'h0; // @[ICache.scala 59:26]
    end else if (5'he == index_addr) begin // @[ICache.scala 114:26]
      if (_block2_T) begin // @[ICache.scala 114:32]
        tag2_14 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 63:28]
        tag2_14 <= tag2_31; // @[ICache.scala 63:28]
      end else begin
        tag2_14 <= _GEN_95;
      end
    end
    if (reset) begin // @[ICache.scala 59:26]
      tag2_15 <= 53'h0; // @[ICache.scala 59:26]
    end else if (5'hf == index_addr) begin // @[ICache.scala 114:26]
      if (_block2_T) begin // @[ICache.scala 114:32]
        tag2_15 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 63:28]
        tag2_15 <= tag2_31; // @[ICache.scala 63:28]
      end else begin
        tag2_15 <= _GEN_95;
      end
    end
    if (reset) begin // @[ICache.scala 59:26]
      tag2_16 <= 53'h0; // @[ICache.scala 59:26]
    end else if (5'h10 == index_addr) begin // @[ICache.scala 114:26]
      if (_block2_T) begin // @[ICache.scala 114:32]
        tag2_16 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 63:28]
        tag2_16 <= tag2_31; // @[ICache.scala 63:28]
      end else begin
        tag2_16 <= _GEN_95;
      end
    end
    if (reset) begin // @[ICache.scala 59:26]
      tag2_17 <= 53'h0; // @[ICache.scala 59:26]
    end else if (5'h11 == index_addr) begin // @[ICache.scala 114:26]
      if (_block2_T) begin // @[ICache.scala 114:32]
        tag2_17 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 63:28]
        tag2_17 <= tag2_31; // @[ICache.scala 63:28]
      end else begin
        tag2_17 <= _GEN_95;
      end
    end
    if (reset) begin // @[ICache.scala 59:26]
      tag2_18 <= 53'h0; // @[ICache.scala 59:26]
    end else if (5'h12 == index_addr) begin // @[ICache.scala 114:26]
      if (_block2_T) begin // @[ICache.scala 114:32]
        tag2_18 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 63:28]
        tag2_18 <= tag2_31; // @[ICache.scala 63:28]
      end else begin
        tag2_18 <= _GEN_95;
      end
    end
    if (reset) begin // @[ICache.scala 59:26]
      tag2_19 <= 53'h0; // @[ICache.scala 59:26]
    end else if (5'h13 == index_addr) begin // @[ICache.scala 114:26]
      if (_block2_T) begin // @[ICache.scala 114:32]
        tag2_19 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 63:28]
        tag2_19 <= tag2_31; // @[ICache.scala 63:28]
      end else begin
        tag2_19 <= _GEN_95;
      end
    end
    if (reset) begin // @[ICache.scala 59:26]
      tag2_20 <= 53'h0; // @[ICache.scala 59:26]
    end else if (5'h14 == index_addr) begin // @[ICache.scala 114:26]
      if (_block2_T) begin // @[ICache.scala 114:32]
        tag2_20 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 63:28]
        tag2_20 <= tag2_31; // @[ICache.scala 63:28]
      end else begin
        tag2_20 <= _GEN_95;
      end
    end
    if (reset) begin // @[ICache.scala 59:26]
      tag2_21 <= 53'h0; // @[ICache.scala 59:26]
    end else if (5'h15 == index_addr) begin // @[ICache.scala 114:26]
      if (_block2_T) begin // @[ICache.scala 114:32]
        tag2_21 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 63:28]
        tag2_21 <= tag2_31; // @[ICache.scala 63:28]
      end else begin
        tag2_21 <= _GEN_95;
      end
    end
    if (reset) begin // @[ICache.scala 59:26]
      tag2_22 <= 53'h0; // @[ICache.scala 59:26]
    end else if (5'h16 == index_addr) begin // @[ICache.scala 114:26]
      if (_block2_T) begin // @[ICache.scala 114:32]
        tag2_22 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 63:28]
        tag2_22 <= tag2_31; // @[ICache.scala 63:28]
      end else begin
        tag2_22 <= _GEN_95;
      end
    end
    if (reset) begin // @[ICache.scala 59:26]
      tag2_23 <= 53'h0; // @[ICache.scala 59:26]
    end else if (5'h17 == index_addr) begin // @[ICache.scala 114:26]
      if (_block2_T) begin // @[ICache.scala 114:32]
        tag2_23 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 63:28]
        tag2_23 <= tag2_31; // @[ICache.scala 63:28]
      end else begin
        tag2_23 <= _GEN_95;
      end
    end
    if (reset) begin // @[ICache.scala 59:26]
      tag2_24 <= 53'h0; // @[ICache.scala 59:26]
    end else if (5'h18 == index_addr) begin // @[ICache.scala 114:26]
      if (_block2_T) begin // @[ICache.scala 114:32]
        tag2_24 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 63:28]
        tag2_24 <= tag2_31; // @[ICache.scala 63:28]
      end else begin
        tag2_24 <= _GEN_95;
      end
    end
    if (reset) begin // @[ICache.scala 59:26]
      tag2_25 <= 53'h0; // @[ICache.scala 59:26]
    end else if (5'h19 == index_addr) begin // @[ICache.scala 114:26]
      if (_block2_T) begin // @[ICache.scala 114:32]
        tag2_25 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 63:28]
        tag2_25 <= tag2_31; // @[ICache.scala 63:28]
      end else begin
        tag2_25 <= _GEN_95;
      end
    end
    if (reset) begin // @[ICache.scala 59:26]
      tag2_26 <= 53'h0; // @[ICache.scala 59:26]
    end else if (5'h1a == index_addr) begin // @[ICache.scala 114:26]
      if (_block2_T) begin // @[ICache.scala 114:32]
        tag2_26 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 63:28]
        tag2_26 <= tag2_31; // @[ICache.scala 63:28]
      end else begin
        tag2_26 <= _GEN_95;
      end
    end
    if (reset) begin // @[ICache.scala 59:26]
      tag2_27 <= 53'h0; // @[ICache.scala 59:26]
    end else if (5'h1b == index_addr) begin // @[ICache.scala 114:26]
      if (_block2_T) begin // @[ICache.scala 114:32]
        tag2_27 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 63:28]
        tag2_27 <= tag2_31; // @[ICache.scala 63:28]
      end else begin
        tag2_27 <= _GEN_95;
      end
    end
    if (reset) begin // @[ICache.scala 59:26]
      tag2_28 <= 53'h0; // @[ICache.scala 59:26]
    end else if (5'h1c == index_addr) begin // @[ICache.scala 114:26]
      if (_block2_T) begin // @[ICache.scala 114:32]
        tag2_28 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 63:28]
        tag2_28 <= tag2_31; // @[ICache.scala 63:28]
      end else begin
        tag2_28 <= _GEN_95;
      end
    end
    if (reset) begin // @[ICache.scala 59:26]
      tag2_29 <= 53'h0; // @[ICache.scala 59:26]
    end else if (5'h1d == index_addr) begin // @[ICache.scala 114:26]
      if (_block2_T) begin // @[ICache.scala 114:32]
        tag2_29 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 63:28]
        tag2_29 <= tag2_31; // @[ICache.scala 63:28]
      end else begin
        tag2_29 <= _GEN_95;
      end
    end
    if (reset) begin // @[ICache.scala 59:26]
      tag2_30 <= 53'h0; // @[ICache.scala 59:26]
    end else if (5'h1e == index_addr) begin // @[ICache.scala 114:26]
      if (_block2_T) begin // @[ICache.scala 114:32]
        tag2_30 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 63:28]
        tag2_30 <= tag2_31; // @[ICache.scala 63:28]
      end else begin
        tag2_30 <= _GEN_95;
      end
    end
    if (reset) begin // @[ICache.scala 59:26]
      tag2_31 <= 53'h0; // @[ICache.scala 59:26]
    end else if (5'h1f == index_addr) begin // @[ICache.scala 114:26]
      if (_block2_T) begin // @[ICache.scala 114:32]
        tag2_31 <= tag_addr;
      end else if (!(5'h1f == index_addr)) begin // @[ICache.scala 63:28]
        tag2_31 <= _GEN_95;
      end
    end
    if (reset) begin // @[ICache.scala 60:26]
      block2_0 <= 512'h0; // @[ICache.scala 60:26]
    end else if (5'h0 == index_addr) begin // @[ICache.scala 113:26]
      if (update & updateway2) begin // @[ICache.scala 113:32]
        block2_0 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 65:39]
        block2_0 <= block2_31; // @[ICache.scala 65:39]
      end else begin
        block2_0 <= _GEN_191;
      end
    end
    if (reset) begin // @[ICache.scala 60:26]
      block2_1 <= 512'h0; // @[ICache.scala 60:26]
    end else if (5'h1 == index_addr) begin // @[ICache.scala 113:26]
      if (update & updateway2) begin // @[ICache.scala 113:32]
        block2_1 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 65:39]
        block2_1 <= block2_31; // @[ICache.scala 65:39]
      end else begin
        block2_1 <= _GEN_191;
      end
    end
    if (reset) begin // @[ICache.scala 60:26]
      block2_2 <= 512'h0; // @[ICache.scala 60:26]
    end else if (5'h2 == index_addr) begin // @[ICache.scala 113:26]
      if (update & updateway2) begin // @[ICache.scala 113:32]
        block2_2 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 65:39]
        block2_2 <= block2_31; // @[ICache.scala 65:39]
      end else begin
        block2_2 <= _GEN_191;
      end
    end
    if (reset) begin // @[ICache.scala 60:26]
      block2_3 <= 512'h0; // @[ICache.scala 60:26]
    end else if (5'h3 == index_addr) begin // @[ICache.scala 113:26]
      if (update & updateway2) begin // @[ICache.scala 113:32]
        block2_3 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 65:39]
        block2_3 <= block2_31; // @[ICache.scala 65:39]
      end else begin
        block2_3 <= _GEN_191;
      end
    end
    if (reset) begin // @[ICache.scala 60:26]
      block2_4 <= 512'h0; // @[ICache.scala 60:26]
    end else if (5'h4 == index_addr) begin // @[ICache.scala 113:26]
      if (update & updateway2) begin // @[ICache.scala 113:32]
        block2_4 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 65:39]
        block2_4 <= block2_31; // @[ICache.scala 65:39]
      end else begin
        block2_4 <= _GEN_191;
      end
    end
    if (reset) begin // @[ICache.scala 60:26]
      block2_5 <= 512'h0; // @[ICache.scala 60:26]
    end else if (5'h5 == index_addr) begin // @[ICache.scala 113:26]
      if (update & updateway2) begin // @[ICache.scala 113:32]
        block2_5 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 65:39]
        block2_5 <= block2_31; // @[ICache.scala 65:39]
      end else begin
        block2_5 <= _GEN_191;
      end
    end
    if (reset) begin // @[ICache.scala 60:26]
      block2_6 <= 512'h0; // @[ICache.scala 60:26]
    end else if (5'h6 == index_addr) begin // @[ICache.scala 113:26]
      if (update & updateway2) begin // @[ICache.scala 113:32]
        block2_6 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 65:39]
        block2_6 <= block2_31; // @[ICache.scala 65:39]
      end else begin
        block2_6 <= _GEN_191;
      end
    end
    if (reset) begin // @[ICache.scala 60:26]
      block2_7 <= 512'h0; // @[ICache.scala 60:26]
    end else if (5'h7 == index_addr) begin // @[ICache.scala 113:26]
      if (update & updateway2) begin // @[ICache.scala 113:32]
        block2_7 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 65:39]
        block2_7 <= block2_31; // @[ICache.scala 65:39]
      end else begin
        block2_7 <= _GEN_191;
      end
    end
    if (reset) begin // @[ICache.scala 60:26]
      block2_8 <= 512'h0; // @[ICache.scala 60:26]
    end else if (5'h8 == index_addr) begin // @[ICache.scala 113:26]
      if (update & updateway2) begin // @[ICache.scala 113:32]
        block2_8 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 65:39]
        block2_8 <= block2_31; // @[ICache.scala 65:39]
      end else begin
        block2_8 <= _GEN_191;
      end
    end
    if (reset) begin // @[ICache.scala 60:26]
      block2_9 <= 512'h0; // @[ICache.scala 60:26]
    end else if (5'h9 == index_addr) begin // @[ICache.scala 113:26]
      if (update & updateway2) begin // @[ICache.scala 113:32]
        block2_9 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 65:39]
        block2_9 <= block2_31; // @[ICache.scala 65:39]
      end else begin
        block2_9 <= _GEN_191;
      end
    end
    if (reset) begin // @[ICache.scala 60:26]
      block2_10 <= 512'h0; // @[ICache.scala 60:26]
    end else if (5'ha == index_addr) begin // @[ICache.scala 113:26]
      if (update & updateway2) begin // @[ICache.scala 113:32]
        block2_10 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 65:39]
        block2_10 <= block2_31; // @[ICache.scala 65:39]
      end else begin
        block2_10 <= _GEN_191;
      end
    end
    if (reset) begin // @[ICache.scala 60:26]
      block2_11 <= 512'h0; // @[ICache.scala 60:26]
    end else if (5'hb == index_addr) begin // @[ICache.scala 113:26]
      if (update & updateway2) begin // @[ICache.scala 113:32]
        block2_11 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 65:39]
        block2_11 <= block2_31; // @[ICache.scala 65:39]
      end else begin
        block2_11 <= _GEN_191;
      end
    end
    if (reset) begin // @[ICache.scala 60:26]
      block2_12 <= 512'h0; // @[ICache.scala 60:26]
    end else if (5'hc == index_addr) begin // @[ICache.scala 113:26]
      if (update & updateway2) begin // @[ICache.scala 113:32]
        block2_12 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 65:39]
        block2_12 <= block2_31; // @[ICache.scala 65:39]
      end else begin
        block2_12 <= _GEN_191;
      end
    end
    if (reset) begin // @[ICache.scala 60:26]
      block2_13 <= 512'h0; // @[ICache.scala 60:26]
    end else if (5'hd == index_addr) begin // @[ICache.scala 113:26]
      if (update & updateway2) begin // @[ICache.scala 113:32]
        block2_13 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 65:39]
        block2_13 <= block2_31; // @[ICache.scala 65:39]
      end else begin
        block2_13 <= _GEN_191;
      end
    end
    if (reset) begin // @[ICache.scala 60:26]
      block2_14 <= 512'h0; // @[ICache.scala 60:26]
    end else if (5'he == index_addr) begin // @[ICache.scala 113:26]
      if (update & updateway2) begin // @[ICache.scala 113:32]
        block2_14 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 65:39]
        block2_14 <= block2_31; // @[ICache.scala 65:39]
      end else begin
        block2_14 <= _GEN_191;
      end
    end
    if (reset) begin // @[ICache.scala 60:26]
      block2_15 <= 512'h0; // @[ICache.scala 60:26]
    end else if (5'hf == index_addr) begin // @[ICache.scala 113:26]
      if (update & updateway2) begin // @[ICache.scala 113:32]
        block2_15 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 65:39]
        block2_15 <= block2_31; // @[ICache.scala 65:39]
      end else begin
        block2_15 <= _GEN_191;
      end
    end
    if (reset) begin // @[ICache.scala 60:26]
      block2_16 <= 512'h0; // @[ICache.scala 60:26]
    end else if (5'h10 == index_addr) begin // @[ICache.scala 113:26]
      if (update & updateway2) begin // @[ICache.scala 113:32]
        block2_16 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 65:39]
        block2_16 <= block2_31; // @[ICache.scala 65:39]
      end else begin
        block2_16 <= _GEN_191;
      end
    end
    if (reset) begin // @[ICache.scala 60:26]
      block2_17 <= 512'h0; // @[ICache.scala 60:26]
    end else if (5'h11 == index_addr) begin // @[ICache.scala 113:26]
      if (update & updateway2) begin // @[ICache.scala 113:32]
        block2_17 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 65:39]
        block2_17 <= block2_31; // @[ICache.scala 65:39]
      end else begin
        block2_17 <= _GEN_191;
      end
    end
    if (reset) begin // @[ICache.scala 60:26]
      block2_18 <= 512'h0; // @[ICache.scala 60:26]
    end else if (5'h12 == index_addr) begin // @[ICache.scala 113:26]
      if (update & updateway2) begin // @[ICache.scala 113:32]
        block2_18 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 65:39]
        block2_18 <= block2_31; // @[ICache.scala 65:39]
      end else begin
        block2_18 <= _GEN_191;
      end
    end
    if (reset) begin // @[ICache.scala 60:26]
      block2_19 <= 512'h0; // @[ICache.scala 60:26]
    end else if (5'h13 == index_addr) begin // @[ICache.scala 113:26]
      if (update & updateway2) begin // @[ICache.scala 113:32]
        block2_19 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 65:39]
        block2_19 <= block2_31; // @[ICache.scala 65:39]
      end else begin
        block2_19 <= _GEN_191;
      end
    end
    if (reset) begin // @[ICache.scala 60:26]
      block2_20 <= 512'h0; // @[ICache.scala 60:26]
    end else if (5'h14 == index_addr) begin // @[ICache.scala 113:26]
      if (update & updateway2) begin // @[ICache.scala 113:32]
        block2_20 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 65:39]
        block2_20 <= block2_31; // @[ICache.scala 65:39]
      end else begin
        block2_20 <= _GEN_191;
      end
    end
    if (reset) begin // @[ICache.scala 60:26]
      block2_21 <= 512'h0; // @[ICache.scala 60:26]
    end else if (5'h15 == index_addr) begin // @[ICache.scala 113:26]
      if (update & updateway2) begin // @[ICache.scala 113:32]
        block2_21 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 65:39]
        block2_21 <= block2_31; // @[ICache.scala 65:39]
      end else begin
        block2_21 <= _GEN_191;
      end
    end
    if (reset) begin // @[ICache.scala 60:26]
      block2_22 <= 512'h0; // @[ICache.scala 60:26]
    end else if (5'h16 == index_addr) begin // @[ICache.scala 113:26]
      if (update & updateway2) begin // @[ICache.scala 113:32]
        block2_22 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 65:39]
        block2_22 <= block2_31; // @[ICache.scala 65:39]
      end else begin
        block2_22 <= _GEN_191;
      end
    end
    if (reset) begin // @[ICache.scala 60:26]
      block2_23 <= 512'h0; // @[ICache.scala 60:26]
    end else if (5'h17 == index_addr) begin // @[ICache.scala 113:26]
      if (update & updateway2) begin // @[ICache.scala 113:32]
        block2_23 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 65:39]
        block2_23 <= block2_31; // @[ICache.scala 65:39]
      end else begin
        block2_23 <= _GEN_191;
      end
    end
    if (reset) begin // @[ICache.scala 60:26]
      block2_24 <= 512'h0; // @[ICache.scala 60:26]
    end else if (5'h18 == index_addr) begin // @[ICache.scala 113:26]
      if (update & updateway2) begin // @[ICache.scala 113:32]
        block2_24 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 65:39]
        block2_24 <= block2_31; // @[ICache.scala 65:39]
      end else begin
        block2_24 <= _GEN_191;
      end
    end
    if (reset) begin // @[ICache.scala 60:26]
      block2_25 <= 512'h0; // @[ICache.scala 60:26]
    end else if (5'h19 == index_addr) begin // @[ICache.scala 113:26]
      if (update & updateway2) begin // @[ICache.scala 113:32]
        block2_25 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 65:39]
        block2_25 <= block2_31; // @[ICache.scala 65:39]
      end else begin
        block2_25 <= _GEN_191;
      end
    end
    if (reset) begin // @[ICache.scala 60:26]
      block2_26 <= 512'h0; // @[ICache.scala 60:26]
    end else if (5'h1a == index_addr) begin // @[ICache.scala 113:26]
      if (update & updateway2) begin // @[ICache.scala 113:32]
        block2_26 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 65:39]
        block2_26 <= block2_31; // @[ICache.scala 65:39]
      end else begin
        block2_26 <= _GEN_191;
      end
    end
    if (reset) begin // @[ICache.scala 60:26]
      block2_27 <= 512'h0; // @[ICache.scala 60:26]
    end else if (5'h1b == index_addr) begin // @[ICache.scala 113:26]
      if (update & updateway2) begin // @[ICache.scala 113:32]
        block2_27 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 65:39]
        block2_27 <= block2_31; // @[ICache.scala 65:39]
      end else begin
        block2_27 <= _GEN_191;
      end
    end
    if (reset) begin // @[ICache.scala 60:26]
      block2_28 <= 512'h0; // @[ICache.scala 60:26]
    end else if (5'h1c == index_addr) begin // @[ICache.scala 113:26]
      if (update & updateway2) begin // @[ICache.scala 113:32]
        block2_28 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 65:39]
        block2_28 <= block2_31; // @[ICache.scala 65:39]
      end else begin
        block2_28 <= _GEN_191;
      end
    end
    if (reset) begin // @[ICache.scala 60:26]
      block2_29 <= 512'h0; // @[ICache.scala 60:26]
    end else if (5'h1d == index_addr) begin // @[ICache.scala 113:26]
      if (update & updateway2) begin // @[ICache.scala 113:32]
        block2_29 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 65:39]
        block2_29 <= block2_31; // @[ICache.scala 65:39]
      end else begin
        block2_29 <= _GEN_191;
      end
    end
    if (reset) begin // @[ICache.scala 60:26]
      block2_30 <= 512'h0; // @[ICache.scala 60:26]
    end else if (5'h1e == index_addr) begin // @[ICache.scala 113:26]
      if (update & updateway2) begin // @[ICache.scala 113:32]
        block2_30 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 65:39]
        block2_30 <= block2_31; // @[ICache.scala 65:39]
      end else begin
        block2_30 <= _GEN_191;
      end
    end
    if (reset) begin // @[ICache.scala 60:26]
      block2_31 <= 512'h0; // @[ICache.scala 60:26]
    end else if (5'h1f == index_addr) begin // @[ICache.scala 113:26]
      if (update & updateway2) begin // @[ICache.scala 113:32]
        block2_31 <= io_axi_data;
      end else if (!(5'h1f == index_addr)) begin // @[ICache.scala 65:39]
        block2_31 <= _GEN_191;
      end
    end
    if (reset) begin // @[ICache.scala 75:24]
      state <= 2'h0; // @[ICache.scala 75:24]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_fence_req) begin // @[ICache.scala 87:31]
        state <= 2'h2; // @[ICache.scala 87:38]
      end else if (~hit & ~not_en_yet) begin // @[ICache.scala 88:43]
        state <= 2'h1; // @[ICache.scala 88:50]
      end
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      if (io_axi_valid) begin // @[ICache.scala 91:32]
        state <= 2'h0; // @[ICache.scala 91:39]
      end
    end else if (_T_5) begin // @[Conditional.scala 39:67]
      state <= _GEN_324;
    end else begin
      state <= _GEN_326;
    end
    not_en_yet <= reset | _not_en_yet_T; // @[ICache.scala 78:30 ICache.scala 78:30 ICache.scala 79:21]
    if (reset) begin // @[ICache.scala 84:28]
      fence_cnt <= 5'h0; // @[ICache.scala 84:28]
    end else if (_T_9 | _T_11) begin // @[ICache.scala 123:59]
      fence_cnt <= _fence_cnt_T_1; // @[ICache.scala 123:70]
    end else begin
      fence_cnt <= 5'h0; // @[ICache.scala 124:26]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  addr = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  v1_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  v1_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  v1_2 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  v1_3 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  v1_4 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  v1_5 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  v1_6 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  v1_7 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  v1_8 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  v1_9 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  v1_10 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  v1_11 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  v1_12 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  v1_13 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  v1_14 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  v1_15 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  v1_16 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  v1_17 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  v1_18 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  v1_19 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  v1_20 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  v1_21 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  v1_22 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  v1_23 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  v1_24 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  v1_25 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  v1_26 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  v1_27 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  v1_28 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  v1_29 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  v1_30 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  v1_31 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  age1_0 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  age1_1 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  age1_2 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  age1_3 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  age1_4 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  age1_5 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  age1_6 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  age1_7 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  age1_8 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  age1_9 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  age1_10 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  age1_11 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  age1_12 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  age1_13 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  age1_14 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  age1_15 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  age1_16 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  age1_17 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  age1_18 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  age1_19 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  age1_20 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  age1_21 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  age1_22 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  age1_23 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  age1_24 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  age1_25 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  age1_26 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  age1_27 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  age1_28 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  age1_29 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  age1_30 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  age1_31 = _RAND_64[0:0];
  _RAND_65 = {2{`RANDOM}};
  tag1_0 = _RAND_65[52:0];
  _RAND_66 = {2{`RANDOM}};
  tag1_1 = _RAND_66[52:0];
  _RAND_67 = {2{`RANDOM}};
  tag1_2 = _RAND_67[52:0];
  _RAND_68 = {2{`RANDOM}};
  tag1_3 = _RAND_68[52:0];
  _RAND_69 = {2{`RANDOM}};
  tag1_4 = _RAND_69[52:0];
  _RAND_70 = {2{`RANDOM}};
  tag1_5 = _RAND_70[52:0];
  _RAND_71 = {2{`RANDOM}};
  tag1_6 = _RAND_71[52:0];
  _RAND_72 = {2{`RANDOM}};
  tag1_7 = _RAND_72[52:0];
  _RAND_73 = {2{`RANDOM}};
  tag1_8 = _RAND_73[52:0];
  _RAND_74 = {2{`RANDOM}};
  tag1_9 = _RAND_74[52:0];
  _RAND_75 = {2{`RANDOM}};
  tag1_10 = _RAND_75[52:0];
  _RAND_76 = {2{`RANDOM}};
  tag1_11 = _RAND_76[52:0];
  _RAND_77 = {2{`RANDOM}};
  tag1_12 = _RAND_77[52:0];
  _RAND_78 = {2{`RANDOM}};
  tag1_13 = _RAND_78[52:0];
  _RAND_79 = {2{`RANDOM}};
  tag1_14 = _RAND_79[52:0];
  _RAND_80 = {2{`RANDOM}};
  tag1_15 = _RAND_80[52:0];
  _RAND_81 = {2{`RANDOM}};
  tag1_16 = _RAND_81[52:0];
  _RAND_82 = {2{`RANDOM}};
  tag1_17 = _RAND_82[52:0];
  _RAND_83 = {2{`RANDOM}};
  tag1_18 = _RAND_83[52:0];
  _RAND_84 = {2{`RANDOM}};
  tag1_19 = _RAND_84[52:0];
  _RAND_85 = {2{`RANDOM}};
  tag1_20 = _RAND_85[52:0];
  _RAND_86 = {2{`RANDOM}};
  tag1_21 = _RAND_86[52:0];
  _RAND_87 = {2{`RANDOM}};
  tag1_22 = _RAND_87[52:0];
  _RAND_88 = {2{`RANDOM}};
  tag1_23 = _RAND_88[52:0];
  _RAND_89 = {2{`RANDOM}};
  tag1_24 = _RAND_89[52:0];
  _RAND_90 = {2{`RANDOM}};
  tag1_25 = _RAND_90[52:0];
  _RAND_91 = {2{`RANDOM}};
  tag1_26 = _RAND_91[52:0];
  _RAND_92 = {2{`RANDOM}};
  tag1_27 = _RAND_92[52:0];
  _RAND_93 = {2{`RANDOM}};
  tag1_28 = _RAND_93[52:0];
  _RAND_94 = {2{`RANDOM}};
  tag1_29 = _RAND_94[52:0];
  _RAND_95 = {2{`RANDOM}};
  tag1_30 = _RAND_95[52:0];
  _RAND_96 = {2{`RANDOM}};
  tag1_31 = _RAND_96[52:0];
  _RAND_97 = {16{`RANDOM}};
  block1_0 = _RAND_97[511:0];
  _RAND_98 = {16{`RANDOM}};
  block1_1 = _RAND_98[511:0];
  _RAND_99 = {16{`RANDOM}};
  block1_2 = _RAND_99[511:0];
  _RAND_100 = {16{`RANDOM}};
  block1_3 = _RAND_100[511:0];
  _RAND_101 = {16{`RANDOM}};
  block1_4 = _RAND_101[511:0];
  _RAND_102 = {16{`RANDOM}};
  block1_5 = _RAND_102[511:0];
  _RAND_103 = {16{`RANDOM}};
  block1_6 = _RAND_103[511:0];
  _RAND_104 = {16{`RANDOM}};
  block1_7 = _RAND_104[511:0];
  _RAND_105 = {16{`RANDOM}};
  block1_8 = _RAND_105[511:0];
  _RAND_106 = {16{`RANDOM}};
  block1_9 = _RAND_106[511:0];
  _RAND_107 = {16{`RANDOM}};
  block1_10 = _RAND_107[511:0];
  _RAND_108 = {16{`RANDOM}};
  block1_11 = _RAND_108[511:0];
  _RAND_109 = {16{`RANDOM}};
  block1_12 = _RAND_109[511:0];
  _RAND_110 = {16{`RANDOM}};
  block1_13 = _RAND_110[511:0];
  _RAND_111 = {16{`RANDOM}};
  block1_14 = _RAND_111[511:0];
  _RAND_112 = {16{`RANDOM}};
  block1_15 = _RAND_112[511:0];
  _RAND_113 = {16{`RANDOM}};
  block1_16 = _RAND_113[511:0];
  _RAND_114 = {16{`RANDOM}};
  block1_17 = _RAND_114[511:0];
  _RAND_115 = {16{`RANDOM}};
  block1_18 = _RAND_115[511:0];
  _RAND_116 = {16{`RANDOM}};
  block1_19 = _RAND_116[511:0];
  _RAND_117 = {16{`RANDOM}};
  block1_20 = _RAND_117[511:0];
  _RAND_118 = {16{`RANDOM}};
  block1_21 = _RAND_118[511:0];
  _RAND_119 = {16{`RANDOM}};
  block1_22 = _RAND_119[511:0];
  _RAND_120 = {16{`RANDOM}};
  block1_23 = _RAND_120[511:0];
  _RAND_121 = {16{`RANDOM}};
  block1_24 = _RAND_121[511:0];
  _RAND_122 = {16{`RANDOM}};
  block1_25 = _RAND_122[511:0];
  _RAND_123 = {16{`RANDOM}};
  block1_26 = _RAND_123[511:0];
  _RAND_124 = {16{`RANDOM}};
  block1_27 = _RAND_124[511:0];
  _RAND_125 = {16{`RANDOM}};
  block1_28 = _RAND_125[511:0];
  _RAND_126 = {16{`RANDOM}};
  block1_29 = _RAND_126[511:0];
  _RAND_127 = {16{`RANDOM}};
  block1_30 = _RAND_127[511:0];
  _RAND_128 = {16{`RANDOM}};
  block1_31 = _RAND_128[511:0];
  _RAND_129 = {1{`RANDOM}};
  v2_0 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  v2_1 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  v2_2 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  v2_3 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  v2_4 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  v2_5 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  v2_6 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  v2_7 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  v2_8 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  v2_9 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  v2_10 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  v2_11 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  v2_12 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  v2_13 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  v2_14 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  v2_15 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  v2_16 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  v2_17 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  v2_18 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  v2_19 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  v2_20 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  v2_21 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  v2_22 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  v2_23 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  v2_24 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  v2_25 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  v2_26 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  v2_27 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  v2_28 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  v2_29 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  v2_30 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  v2_31 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  age2_0 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  age2_1 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  age2_2 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  age2_3 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  age2_4 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  age2_5 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  age2_6 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  age2_7 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  age2_8 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  age2_9 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  age2_10 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  age2_11 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  age2_12 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  age2_13 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  age2_14 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  age2_15 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  age2_16 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  age2_17 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  age2_18 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  age2_19 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  age2_20 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  age2_21 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  age2_22 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  age2_23 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  age2_24 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  age2_25 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  age2_26 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  age2_27 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  age2_28 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  age2_29 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  age2_30 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  age2_31 = _RAND_192[0:0];
  _RAND_193 = {2{`RANDOM}};
  tag2_0 = _RAND_193[52:0];
  _RAND_194 = {2{`RANDOM}};
  tag2_1 = _RAND_194[52:0];
  _RAND_195 = {2{`RANDOM}};
  tag2_2 = _RAND_195[52:0];
  _RAND_196 = {2{`RANDOM}};
  tag2_3 = _RAND_196[52:0];
  _RAND_197 = {2{`RANDOM}};
  tag2_4 = _RAND_197[52:0];
  _RAND_198 = {2{`RANDOM}};
  tag2_5 = _RAND_198[52:0];
  _RAND_199 = {2{`RANDOM}};
  tag2_6 = _RAND_199[52:0];
  _RAND_200 = {2{`RANDOM}};
  tag2_7 = _RAND_200[52:0];
  _RAND_201 = {2{`RANDOM}};
  tag2_8 = _RAND_201[52:0];
  _RAND_202 = {2{`RANDOM}};
  tag2_9 = _RAND_202[52:0];
  _RAND_203 = {2{`RANDOM}};
  tag2_10 = _RAND_203[52:0];
  _RAND_204 = {2{`RANDOM}};
  tag2_11 = _RAND_204[52:0];
  _RAND_205 = {2{`RANDOM}};
  tag2_12 = _RAND_205[52:0];
  _RAND_206 = {2{`RANDOM}};
  tag2_13 = _RAND_206[52:0];
  _RAND_207 = {2{`RANDOM}};
  tag2_14 = _RAND_207[52:0];
  _RAND_208 = {2{`RANDOM}};
  tag2_15 = _RAND_208[52:0];
  _RAND_209 = {2{`RANDOM}};
  tag2_16 = _RAND_209[52:0];
  _RAND_210 = {2{`RANDOM}};
  tag2_17 = _RAND_210[52:0];
  _RAND_211 = {2{`RANDOM}};
  tag2_18 = _RAND_211[52:0];
  _RAND_212 = {2{`RANDOM}};
  tag2_19 = _RAND_212[52:0];
  _RAND_213 = {2{`RANDOM}};
  tag2_20 = _RAND_213[52:0];
  _RAND_214 = {2{`RANDOM}};
  tag2_21 = _RAND_214[52:0];
  _RAND_215 = {2{`RANDOM}};
  tag2_22 = _RAND_215[52:0];
  _RAND_216 = {2{`RANDOM}};
  tag2_23 = _RAND_216[52:0];
  _RAND_217 = {2{`RANDOM}};
  tag2_24 = _RAND_217[52:0];
  _RAND_218 = {2{`RANDOM}};
  tag2_25 = _RAND_218[52:0];
  _RAND_219 = {2{`RANDOM}};
  tag2_26 = _RAND_219[52:0];
  _RAND_220 = {2{`RANDOM}};
  tag2_27 = _RAND_220[52:0];
  _RAND_221 = {2{`RANDOM}};
  tag2_28 = _RAND_221[52:0];
  _RAND_222 = {2{`RANDOM}};
  tag2_29 = _RAND_222[52:0];
  _RAND_223 = {2{`RANDOM}};
  tag2_30 = _RAND_223[52:0];
  _RAND_224 = {2{`RANDOM}};
  tag2_31 = _RAND_224[52:0];
  _RAND_225 = {16{`RANDOM}};
  block2_0 = _RAND_225[511:0];
  _RAND_226 = {16{`RANDOM}};
  block2_1 = _RAND_226[511:0];
  _RAND_227 = {16{`RANDOM}};
  block2_2 = _RAND_227[511:0];
  _RAND_228 = {16{`RANDOM}};
  block2_3 = _RAND_228[511:0];
  _RAND_229 = {16{`RANDOM}};
  block2_4 = _RAND_229[511:0];
  _RAND_230 = {16{`RANDOM}};
  block2_5 = _RAND_230[511:0];
  _RAND_231 = {16{`RANDOM}};
  block2_6 = _RAND_231[511:0];
  _RAND_232 = {16{`RANDOM}};
  block2_7 = _RAND_232[511:0];
  _RAND_233 = {16{`RANDOM}};
  block2_8 = _RAND_233[511:0];
  _RAND_234 = {16{`RANDOM}};
  block2_9 = _RAND_234[511:0];
  _RAND_235 = {16{`RANDOM}};
  block2_10 = _RAND_235[511:0];
  _RAND_236 = {16{`RANDOM}};
  block2_11 = _RAND_236[511:0];
  _RAND_237 = {16{`RANDOM}};
  block2_12 = _RAND_237[511:0];
  _RAND_238 = {16{`RANDOM}};
  block2_13 = _RAND_238[511:0];
  _RAND_239 = {16{`RANDOM}};
  block2_14 = _RAND_239[511:0];
  _RAND_240 = {16{`RANDOM}};
  block2_15 = _RAND_240[511:0];
  _RAND_241 = {16{`RANDOM}};
  block2_16 = _RAND_241[511:0];
  _RAND_242 = {16{`RANDOM}};
  block2_17 = _RAND_242[511:0];
  _RAND_243 = {16{`RANDOM}};
  block2_18 = _RAND_243[511:0];
  _RAND_244 = {16{`RANDOM}};
  block2_19 = _RAND_244[511:0];
  _RAND_245 = {16{`RANDOM}};
  block2_20 = _RAND_245[511:0];
  _RAND_246 = {16{`RANDOM}};
  block2_21 = _RAND_246[511:0];
  _RAND_247 = {16{`RANDOM}};
  block2_22 = _RAND_247[511:0];
  _RAND_248 = {16{`RANDOM}};
  block2_23 = _RAND_248[511:0];
  _RAND_249 = {16{`RANDOM}};
  block2_24 = _RAND_249[511:0];
  _RAND_250 = {16{`RANDOM}};
  block2_25 = _RAND_250[511:0];
  _RAND_251 = {16{`RANDOM}};
  block2_26 = _RAND_251[511:0];
  _RAND_252 = {16{`RANDOM}};
  block2_27 = _RAND_252[511:0];
  _RAND_253 = {16{`RANDOM}};
  block2_28 = _RAND_253[511:0];
  _RAND_254 = {16{`RANDOM}};
  block2_29 = _RAND_254[511:0];
  _RAND_255 = {16{`RANDOM}};
  block2_30 = _RAND_255[511:0];
  _RAND_256 = {16{`RANDOM}};
  block2_31 = _RAND_256[511:0];
  _RAND_257 = {1{`RANDOM}};
  state = _RAND_257[1:0];
  _RAND_258 = {1{`RANDOM}};
  not_en_yet = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  fence_cnt = _RAND_259[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DCache(
  input          clock,
  input          reset,
  input          io_dmem_en,
  input          io_dmem_op,
  input  [63:0]  io_dmem_addr,
  input  [63:0]  io_dmem_wdata,
  input  [7:0]   io_dmem_wmask,
  output         io_dmem_ok,
  output [63:0]  io_dmem_rdata,
  output         io_axi_req,
  output [63:0]  io_axi_raddr,
  input          io_axi_rvalid,
  input  [511:0] io_axi_rdata,
  output         io_axi_weq,
  output [63:0]  io_axi_waddr,
  output [511:0] io_axi_wdata,
  input          io_axi_wdone,
  input          io_fence_req,
  output         io_fence_done
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [63:0] _RAND_100;
  reg [63:0] _RAND_101;
  reg [63:0] _RAND_102;
  reg [63:0] _RAND_103;
  reg [63:0] _RAND_104;
  reg [63:0] _RAND_105;
  reg [63:0] _RAND_106;
  reg [63:0] _RAND_107;
  reg [63:0] _RAND_108;
  reg [63:0] _RAND_109;
  reg [63:0] _RAND_110;
  reg [63:0] _RAND_111;
  reg [63:0] _RAND_112;
  reg [63:0] _RAND_113;
  reg [63:0] _RAND_114;
  reg [63:0] _RAND_115;
  reg [63:0] _RAND_116;
  reg [63:0] _RAND_117;
  reg [63:0] _RAND_118;
  reg [63:0] _RAND_119;
  reg [63:0] _RAND_120;
  reg [63:0] _RAND_121;
  reg [63:0] _RAND_122;
  reg [63:0] _RAND_123;
  reg [63:0] _RAND_124;
  reg [63:0] _RAND_125;
  reg [63:0] _RAND_126;
  reg [63:0] _RAND_127;
  reg [63:0] _RAND_128;
  reg [63:0] _RAND_129;
  reg [63:0] _RAND_130;
  reg [63:0] _RAND_131;
  reg [511:0] _RAND_132;
  reg [511:0] _RAND_133;
  reg [511:0] _RAND_134;
  reg [511:0] _RAND_135;
  reg [511:0] _RAND_136;
  reg [511:0] _RAND_137;
  reg [511:0] _RAND_138;
  reg [511:0] _RAND_139;
  reg [511:0] _RAND_140;
  reg [511:0] _RAND_141;
  reg [511:0] _RAND_142;
  reg [511:0] _RAND_143;
  reg [511:0] _RAND_144;
  reg [511:0] _RAND_145;
  reg [511:0] _RAND_146;
  reg [511:0] _RAND_147;
  reg [511:0] _RAND_148;
  reg [511:0] _RAND_149;
  reg [511:0] _RAND_150;
  reg [511:0] _RAND_151;
  reg [511:0] _RAND_152;
  reg [511:0] _RAND_153;
  reg [511:0] _RAND_154;
  reg [511:0] _RAND_155;
  reg [511:0] _RAND_156;
  reg [511:0] _RAND_157;
  reg [511:0] _RAND_158;
  reg [511:0] _RAND_159;
  reg [511:0] _RAND_160;
  reg [511:0] _RAND_161;
  reg [511:0] _RAND_162;
  reg [511:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [63:0] _RAND_260;
  reg [63:0] _RAND_261;
  reg [63:0] _RAND_262;
  reg [63:0] _RAND_263;
  reg [63:0] _RAND_264;
  reg [63:0] _RAND_265;
  reg [63:0] _RAND_266;
  reg [63:0] _RAND_267;
  reg [63:0] _RAND_268;
  reg [63:0] _RAND_269;
  reg [63:0] _RAND_270;
  reg [63:0] _RAND_271;
  reg [63:0] _RAND_272;
  reg [63:0] _RAND_273;
  reg [63:0] _RAND_274;
  reg [63:0] _RAND_275;
  reg [63:0] _RAND_276;
  reg [63:0] _RAND_277;
  reg [63:0] _RAND_278;
  reg [63:0] _RAND_279;
  reg [63:0] _RAND_280;
  reg [63:0] _RAND_281;
  reg [63:0] _RAND_282;
  reg [63:0] _RAND_283;
  reg [63:0] _RAND_284;
  reg [63:0] _RAND_285;
  reg [63:0] _RAND_286;
  reg [63:0] _RAND_287;
  reg [63:0] _RAND_288;
  reg [63:0] _RAND_289;
  reg [63:0] _RAND_290;
  reg [63:0] _RAND_291;
  reg [511:0] _RAND_292;
  reg [511:0] _RAND_293;
  reg [511:0] _RAND_294;
  reg [511:0] _RAND_295;
  reg [511:0] _RAND_296;
  reg [511:0] _RAND_297;
  reg [511:0] _RAND_298;
  reg [511:0] _RAND_299;
  reg [511:0] _RAND_300;
  reg [511:0] _RAND_301;
  reg [511:0] _RAND_302;
  reg [511:0] _RAND_303;
  reg [511:0] _RAND_304;
  reg [511:0] _RAND_305;
  reg [511:0] _RAND_306;
  reg [511:0] _RAND_307;
  reg [511:0] _RAND_308;
  reg [511:0] _RAND_309;
  reg [511:0] _RAND_310;
  reg [511:0] _RAND_311;
  reg [511:0] _RAND_312;
  reg [511:0] _RAND_313;
  reg [511:0] _RAND_314;
  reg [511:0] _RAND_315;
  reg [511:0] _RAND_316;
  reg [511:0] _RAND_317;
  reg [511:0] _RAND_318;
  reg [511:0] _RAND_319;
  reg [511:0] _RAND_320;
  reg [511:0] _RAND_321;
  reg [511:0] _RAND_322;
  reg [511:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
`endif // RANDOMIZE_REG_INIT
  wire  _op_T = io_dmem_en & io_dmem_ok; // @[DCache.scala 42:66]
  reg  op; // @[Reg.scala 27:20]
  wire [63:0] _addr_T = io_dmem_addr & 64'hfffffffffffffff8; // @[DCache.scala 43:42]
  reg [63:0] addr; // @[Reg.scala 27:20]
  reg [63:0] wdata; // @[Reg.scala 27:20]
  reg [7:0] wm; // @[Reg.scala 27:20]
  wire [52:0] tag_addr = addr[63:11]; // @[DCache.scala 48:27]
  wire [4:0] index_addr = addr[10:6]; // @[DCache.scala 49:27]
  wire [5:0] offset_addr = addr[5:0]; // @[DCache.scala 50:27]
  reg  v1_0; // @[DCache.scala 52:26]
  reg  v1_1; // @[DCache.scala 52:26]
  reg  v1_2; // @[DCache.scala 52:26]
  reg  v1_3; // @[DCache.scala 52:26]
  reg  v1_4; // @[DCache.scala 52:26]
  reg  v1_5; // @[DCache.scala 52:26]
  reg  v1_6; // @[DCache.scala 52:26]
  reg  v1_7; // @[DCache.scala 52:26]
  reg  v1_8; // @[DCache.scala 52:26]
  reg  v1_9; // @[DCache.scala 52:26]
  reg  v1_10; // @[DCache.scala 52:26]
  reg  v1_11; // @[DCache.scala 52:26]
  reg  v1_12; // @[DCache.scala 52:26]
  reg  v1_13; // @[DCache.scala 52:26]
  reg  v1_14; // @[DCache.scala 52:26]
  reg  v1_15; // @[DCache.scala 52:26]
  reg  v1_16; // @[DCache.scala 52:26]
  reg  v1_17; // @[DCache.scala 52:26]
  reg  v1_18; // @[DCache.scala 52:26]
  reg  v1_19; // @[DCache.scala 52:26]
  reg  v1_20; // @[DCache.scala 52:26]
  reg  v1_21; // @[DCache.scala 52:26]
  reg  v1_22; // @[DCache.scala 52:26]
  reg  v1_23; // @[DCache.scala 52:26]
  reg  v1_24; // @[DCache.scala 52:26]
  reg  v1_25; // @[DCache.scala 52:26]
  reg  v1_26; // @[DCache.scala 52:26]
  reg  v1_27; // @[DCache.scala 52:26]
  reg  v1_28; // @[DCache.scala 52:26]
  reg  v1_29; // @[DCache.scala 52:26]
  reg  v1_30; // @[DCache.scala 52:26]
  reg  v1_31; // @[DCache.scala 52:26]
  reg  d1_0; // @[DCache.scala 53:26]
  reg  d1_1; // @[DCache.scala 53:26]
  reg  d1_2; // @[DCache.scala 53:26]
  reg  d1_3; // @[DCache.scala 53:26]
  reg  d1_4; // @[DCache.scala 53:26]
  reg  d1_5; // @[DCache.scala 53:26]
  reg  d1_6; // @[DCache.scala 53:26]
  reg  d1_7; // @[DCache.scala 53:26]
  reg  d1_8; // @[DCache.scala 53:26]
  reg  d1_9; // @[DCache.scala 53:26]
  reg  d1_10; // @[DCache.scala 53:26]
  reg  d1_11; // @[DCache.scala 53:26]
  reg  d1_12; // @[DCache.scala 53:26]
  reg  d1_13; // @[DCache.scala 53:26]
  reg  d1_14; // @[DCache.scala 53:26]
  reg  d1_15; // @[DCache.scala 53:26]
  reg  d1_16; // @[DCache.scala 53:26]
  reg  d1_17; // @[DCache.scala 53:26]
  reg  d1_18; // @[DCache.scala 53:26]
  reg  d1_19; // @[DCache.scala 53:26]
  reg  d1_20; // @[DCache.scala 53:26]
  reg  d1_21; // @[DCache.scala 53:26]
  reg  d1_22; // @[DCache.scala 53:26]
  reg  d1_23; // @[DCache.scala 53:26]
  reg  d1_24; // @[DCache.scala 53:26]
  reg  d1_25; // @[DCache.scala 53:26]
  reg  d1_26; // @[DCache.scala 53:26]
  reg  d1_27; // @[DCache.scala 53:26]
  reg  d1_28; // @[DCache.scala 53:26]
  reg  d1_29; // @[DCache.scala 53:26]
  reg  d1_30; // @[DCache.scala 53:26]
  reg  d1_31; // @[DCache.scala 53:26]
  reg  age1_0; // @[DCache.scala 54:26]
  reg  age1_1; // @[DCache.scala 54:26]
  reg  age1_2; // @[DCache.scala 54:26]
  reg  age1_3; // @[DCache.scala 54:26]
  reg  age1_4; // @[DCache.scala 54:26]
  reg  age1_5; // @[DCache.scala 54:26]
  reg  age1_6; // @[DCache.scala 54:26]
  reg  age1_7; // @[DCache.scala 54:26]
  reg  age1_8; // @[DCache.scala 54:26]
  reg  age1_9; // @[DCache.scala 54:26]
  reg  age1_10; // @[DCache.scala 54:26]
  reg  age1_11; // @[DCache.scala 54:26]
  reg  age1_12; // @[DCache.scala 54:26]
  reg  age1_13; // @[DCache.scala 54:26]
  reg  age1_14; // @[DCache.scala 54:26]
  reg  age1_15; // @[DCache.scala 54:26]
  reg  age1_16; // @[DCache.scala 54:26]
  reg  age1_17; // @[DCache.scala 54:26]
  reg  age1_18; // @[DCache.scala 54:26]
  reg  age1_19; // @[DCache.scala 54:26]
  reg  age1_20; // @[DCache.scala 54:26]
  reg  age1_21; // @[DCache.scala 54:26]
  reg  age1_22; // @[DCache.scala 54:26]
  reg  age1_23; // @[DCache.scala 54:26]
  reg  age1_24; // @[DCache.scala 54:26]
  reg  age1_25; // @[DCache.scala 54:26]
  reg  age1_26; // @[DCache.scala 54:26]
  reg  age1_27; // @[DCache.scala 54:26]
  reg  age1_28; // @[DCache.scala 54:26]
  reg  age1_29; // @[DCache.scala 54:26]
  reg  age1_30; // @[DCache.scala 54:26]
  reg  age1_31; // @[DCache.scala 54:26]
  reg [52:0] tag1_0; // @[DCache.scala 55:26]
  reg [52:0] tag1_1; // @[DCache.scala 55:26]
  reg [52:0] tag1_2; // @[DCache.scala 55:26]
  reg [52:0] tag1_3; // @[DCache.scala 55:26]
  reg [52:0] tag1_4; // @[DCache.scala 55:26]
  reg [52:0] tag1_5; // @[DCache.scala 55:26]
  reg [52:0] tag1_6; // @[DCache.scala 55:26]
  reg [52:0] tag1_7; // @[DCache.scala 55:26]
  reg [52:0] tag1_8; // @[DCache.scala 55:26]
  reg [52:0] tag1_9; // @[DCache.scala 55:26]
  reg [52:0] tag1_10; // @[DCache.scala 55:26]
  reg [52:0] tag1_11; // @[DCache.scala 55:26]
  reg [52:0] tag1_12; // @[DCache.scala 55:26]
  reg [52:0] tag1_13; // @[DCache.scala 55:26]
  reg [52:0] tag1_14; // @[DCache.scala 55:26]
  reg [52:0] tag1_15; // @[DCache.scala 55:26]
  reg [52:0] tag1_16; // @[DCache.scala 55:26]
  reg [52:0] tag1_17; // @[DCache.scala 55:26]
  reg [52:0] tag1_18; // @[DCache.scala 55:26]
  reg [52:0] tag1_19; // @[DCache.scala 55:26]
  reg [52:0] tag1_20; // @[DCache.scala 55:26]
  reg [52:0] tag1_21; // @[DCache.scala 55:26]
  reg [52:0] tag1_22; // @[DCache.scala 55:26]
  reg [52:0] tag1_23; // @[DCache.scala 55:26]
  reg [52:0] tag1_24; // @[DCache.scala 55:26]
  reg [52:0] tag1_25; // @[DCache.scala 55:26]
  reg [52:0] tag1_26; // @[DCache.scala 55:26]
  reg [52:0] tag1_27; // @[DCache.scala 55:26]
  reg [52:0] tag1_28; // @[DCache.scala 55:26]
  reg [52:0] tag1_29; // @[DCache.scala 55:26]
  reg [52:0] tag1_30; // @[DCache.scala 55:26]
  reg [52:0] tag1_31; // @[DCache.scala 55:26]
  reg [511:0] block1_0; // @[DCache.scala 56:26]
  reg [511:0] block1_1; // @[DCache.scala 56:26]
  reg [511:0] block1_2; // @[DCache.scala 56:26]
  reg [511:0] block1_3; // @[DCache.scala 56:26]
  reg [511:0] block1_4; // @[DCache.scala 56:26]
  reg [511:0] block1_5; // @[DCache.scala 56:26]
  reg [511:0] block1_6; // @[DCache.scala 56:26]
  reg [511:0] block1_7; // @[DCache.scala 56:26]
  reg [511:0] block1_8; // @[DCache.scala 56:26]
  reg [511:0] block1_9; // @[DCache.scala 56:26]
  reg [511:0] block1_10; // @[DCache.scala 56:26]
  reg [511:0] block1_11; // @[DCache.scala 56:26]
  reg [511:0] block1_12; // @[DCache.scala 56:26]
  reg [511:0] block1_13; // @[DCache.scala 56:26]
  reg [511:0] block1_14; // @[DCache.scala 56:26]
  reg [511:0] block1_15; // @[DCache.scala 56:26]
  reg [511:0] block1_16; // @[DCache.scala 56:26]
  reg [511:0] block1_17; // @[DCache.scala 56:26]
  reg [511:0] block1_18; // @[DCache.scala 56:26]
  reg [511:0] block1_19; // @[DCache.scala 56:26]
  reg [511:0] block1_20; // @[DCache.scala 56:26]
  reg [511:0] block1_21; // @[DCache.scala 56:26]
  reg [511:0] block1_22; // @[DCache.scala 56:26]
  reg [511:0] block1_23; // @[DCache.scala 56:26]
  reg [511:0] block1_24; // @[DCache.scala 56:26]
  reg [511:0] block1_25; // @[DCache.scala 56:26]
  reg [511:0] block1_26; // @[DCache.scala 56:26]
  reg [511:0] block1_27; // @[DCache.scala 56:26]
  reg [511:0] block1_28; // @[DCache.scala 56:26]
  reg [511:0] block1_29; // @[DCache.scala 56:26]
  reg [511:0] block1_30; // @[DCache.scala 56:26]
  reg [511:0] block1_31; // @[DCache.scala 56:26]
  reg  v2_0; // @[DCache.scala 57:26]
  reg  v2_1; // @[DCache.scala 57:26]
  reg  v2_2; // @[DCache.scala 57:26]
  reg  v2_3; // @[DCache.scala 57:26]
  reg  v2_4; // @[DCache.scala 57:26]
  reg  v2_5; // @[DCache.scala 57:26]
  reg  v2_6; // @[DCache.scala 57:26]
  reg  v2_7; // @[DCache.scala 57:26]
  reg  v2_8; // @[DCache.scala 57:26]
  reg  v2_9; // @[DCache.scala 57:26]
  reg  v2_10; // @[DCache.scala 57:26]
  reg  v2_11; // @[DCache.scala 57:26]
  reg  v2_12; // @[DCache.scala 57:26]
  reg  v2_13; // @[DCache.scala 57:26]
  reg  v2_14; // @[DCache.scala 57:26]
  reg  v2_15; // @[DCache.scala 57:26]
  reg  v2_16; // @[DCache.scala 57:26]
  reg  v2_17; // @[DCache.scala 57:26]
  reg  v2_18; // @[DCache.scala 57:26]
  reg  v2_19; // @[DCache.scala 57:26]
  reg  v2_20; // @[DCache.scala 57:26]
  reg  v2_21; // @[DCache.scala 57:26]
  reg  v2_22; // @[DCache.scala 57:26]
  reg  v2_23; // @[DCache.scala 57:26]
  reg  v2_24; // @[DCache.scala 57:26]
  reg  v2_25; // @[DCache.scala 57:26]
  reg  v2_26; // @[DCache.scala 57:26]
  reg  v2_27; // @[DCache.scala 57:26]
  reg  v2_28; // @[DCache.scala 57:26]
  reg  v2_29; // @[DCache.scala 57:26]
  reg  v2_30; // @[DCache.scala 57:26]
  reg  v2_31; // @[DCache.scala 57:26]
  reg  d2_0; // @[DCache.scala 58:26]
  reg  d2_1; // @[DCache.scala 58:26]
  reg  d2_2; // @[DCache.scala 58:26]
  reg  d2_3; // @[DCache.scala 58:26]
  reg  d2_4; // @[DCache.scala 58:26]
  reg  d2_5; // @[DCache.scala 58:26]
  reg  d2_6; // @[DCache.scala 58:26]
  reg  d2_7; // @[DCache.scala 58:26]
  reg  d2_8; // @[DCache.scala 58:26]
  reg  d2_9; // @[DCache.scala 58:26]
  reg  d2_10; // @[DCache.scala 58:26]
  reg  d2_11; // @[DCache.scala 58:26]
  reg  d2_12; // @[DCache.scala 58:26]
  reg  d2_13; // @[DCache.scala 58:26]
  reg  d2_14; // @[DCache.scala 58:26]
  reg  d2_15; // @[DCache.scala 58:26]
  reg  d2_16; // @[DCache.scala 58:26]
  reg  d2_17; // @[DCache.scala 58:26]
  reg  d2_18; // @[DCache.scala 58:26]
  reg  d2_19; // @[DCache.scala 58:26]
  reg  d2_20; // @[DCache.scala 58:26]
  reg  d2_21; // @[DCache.scala 58:26]
  reg  d2_22; // @[DCache.scala 58:26]
  reg  d2_23; // @[DCache.scala 58:26]
  reg  d2_24; // @[DCache.scala 58:26]
  reg  d2_25; // @[DCache.scala 58:26]
  reg  d2_26; // @[DCache.scala 58:26]
  reg  d2_27; // @[DCache.scala 58:26]
  reg  d2_28; // @[DCache.scala 58:26]
  reg  d2_29; // @[DCache.scala 58:26]
  reg  d2_30; // @[DCache.scala 58:26]
  reg  d2_31; // @[DCache.scala 58:26]
  reg  age2_0; // @[DCache.scala 59:26]
  reg  age2_1; // @[DCache.scala 59:26]
  reg  age2_2; // @[DCache.scala 59:26]
  reg  age2_3; // @[DCache.scala 59:26]
  reg  age2_4; // @[DCache.scala 59:26]
  reg  age2_5; // @[DCache.scala 59:26]
  reg  age2_6; // @[DCache.scala 59:26]
  reg  age2_7; // @[DCache.scala 59:26]
  reg  age2_8; // @[DCache.scala 59:26]
  reg  age2_9; // @[DCache.scala 59:26]
  reg  age2_10; // @[DCache.scala 59:26]
  reg  age2_11; // @[DCache.scala 59:26]
  reg  age2_12; // @[DCache.scala 59:26]
  reg  age2_13; // @[DCache.scala 59:26]
  reg  age2_14; // @[DCache.scala 59:26]
  reg  age2_15; // @[DCache.scala 59:26]
  reg  age2_16; // @[DCache.scala 59:26]
  reg  age2_17; // @[DCache.scala 59:26]
  reg  age2_18; // @[DCache.scala 59:26]
  reg  age2_19; // @[DCache.scala 59:26]
  reg  age2_20; // @[DCache.scala 59:26]
  reg  age2_21; // @[DCache.scala 59:26]
  reg  age2_22; // @[DCache.scala 59:26]
  reg  age2_23; // @[DCache.scala 59:26]
  reg  age2_24; // @[DCache.scala 59:26]
  reg  age2_25; // @[DCache.scala 59:26]
  reg  age2_26; // @[DCache.scala 59:26]
  reg  age2_27; // @[DCache.scala 59:26]
  reg  age2_28; // @[DCache.scala 59:26]
  reg  age2_29; // @[DCache.scala 59:26]
  reg  age2_30; // @[DCache.scala 59:26]
  reg  age2_31; // @[DCache.scala 59:26]
  reg [52:0] tag2_0; // @[DCache.scala 60:26]
  reg [52:0] tag2_1; // @[DCache.scala 60:26]
  reg [52:0] tag2_2; // @[DCache.scala 60:26]
  reg [52:0] tag2_3; // @[DCache.scala 60:26]
  reg [52:0] tag2_4; // @[DCache.scala 60:26]
  reg [52:0] tag2_5; // @[DCache.scala 60:26]
  reg [52:0] tag2_6; // @[DCache.scala 60:26]
  reg [52:0] tag2_7; // @[DCache.scala 60:26]
  reg [52:0] tag2_8; // @[DCache.scala 60:26]
  reg [52:0] tag2_9; // @[DCache.scala 60:26]
  reg [52:0] tag2_10; // @[DCache.scala 60:26]
  reg [52:0] tag2_11; // @[DCache.scala 60:26]
  reg [52:0] tag2_12; // @[DCache.scala 60:26]
  reg [52:0] tag2_13; // @[DCache.scala 60:26]
  reg [52:0] tag2_14; // @[DCache.scala 60:26]
  reg [52:0] tag2_15; // @[DCache.scala 60:26]
  reg [52:0] tag2_16; // @[DCache.scala 60:26]
  reg [52:0] tag2_17; // @[DCache.scala 60:26]
  reg [52:0] tag2_18; // @[DCache.scala 60:26]
  reg [52:0] tag2_19; // @[DCache.scala 60:26]
  reg [52:0] tag2_20; // @[DCache.scala 60:26]
  reg [52:0] tag2_21; // @[DCache.scala 60:26]
  reg [52:0] tag2_22; // @[DCache.scala 60:26]
  reg [52:0] tag2_23; // @[DCache.scala 60:26]
  reg [52:0] tag2_24; // @[DCache.scala 60:26]
  reg [52:0] tag2_25; // @[DCache.scala 60:26]
  reg [52:0] tag2_26; // @[DCache.scala 60:26]
  reg [52:0] tag2_27; // @[DCache.scala 60:26]
  reg [52:0] tag2_28; // @[DCache.scala 60:26]
  reg [52:0] tag2_29; // @[DCache.scala 60:26]
  reg [52:0] tag2_30; // @[DCache.scala 60:26]
  reg [52:0] tag2_31; // @[DCache.scala 60:26]
  reg [511:0] block2_0; // @[DCache.scala 61:26]
  reg [511:0] block2_1; // @[DCache.scala 61:26]
  reg [511:0] block2_2; // @[DCache.scala 61:26]
  reg [511:0] block2_3; // @[DCache.scala 61:26]
  reg [511:0] block2_4; // @[DCache.scala 61:26]
  reg [511:0] block2_5; // @[DCache.scala 61:26]
  reg [511:0] block2_6; // @[DCache.scala 61:26]
  reg [511:0] block2_7; // @[DCache.scala 61:26]
  reg [511:0] block2_8; // @[DCache.scala 61:26]
  reg [511:0] block2_9; // @[DCache.scala 61:26]
  reg [511:0] block2_10; // @[DCache.scala 61:26]
  reg [511:0] block2_11; // @[DCache.scala 61:26]
  reg [511:0] block2_12; // @[DCache.scala 61:26]
  reg [511:0] block2_13; // @[DCache.scala 61:26]
  reg [511:0] block2_14; // @[DCache.scala 61:26]
  reg [511:0] block2_15; // @[DCache.scala 61:26]
  reg [511:0] block2_16; // @[DCache.scala 61:26]
  reg [511:0] block2_17; // @[DCache.scala 61:26]
  reg [511:0] block2_18; // @[DCache.scala 61:26]
  reg [511:0] block2_19; // @[DCache.scala 61:26]
  reg [511:0] block2_20; // @[DCache.scala 61:26]
  reg [511:0] block2_21; // @[DCache.scala 61:26]
  reg [511:0] block2_22; // @[DCache.scala 61:26]
  reg [511:0] block2_23; // @[DCache.scala 61:26]
  reg [511:0] block2_24; // @[DCache.scala 61:26]
  reg [511:0] block2_25; // @[DCache.scala 61:26]
  reg [511:0] block2_26; // @[DCache.scala 61:26]
  reg [511:0] block2_27; // @[DCache.scala 61:26]
  reg [511:0] block2_28; // @[DCache.scala 61:26]
  reg [511:0] block2_29; // @[DCache.scala 61:26]
  reg [511:0] block2_30; // @[DCache.scala 61:26]
  reg [511:0] block2_31; // @[DCache.scala 61:26]
  wire [52:0] _GEN_5 = 5'h1 == index_addr ? tag1_1 : tag1_0; // @[DCache.scala 63:28 DCache.scala 63:28]
  wire [52:0] _GEN_6 = 5'h2 == index_addr ? tag1_2 : _GEN_5; // @[DCache.scala 63:28 DCache.scala 63:28]
  wire [52:0] _GEN_7 = 5'h3 == index_addr ? tag1_3 : _GEN_6; // @[DCache.scala 63:28 DCache.scala 63:28]
  wire [52:0] _GEN_8 = 5'h4 == index_addr ? tag1_4 : _GEN_7; // @[DCache.scala 63:28 DCache.scala 63:28]
  wire [52:0] _GEN_9 = 5'h5 == index_addr ? tag1_5 : _GEN_8; // @[DCache.scala 63:28 DCache.scala 63:28]
  wire [52:0] _GEN_10 = 5'h6 == index_addr ? tag1_6 : _GEN_9; // @[DCache.scala 63:28 DCache.scala 63:28]
  wire [52:0] _GEN_11 = 5'h7 == index_addr ? tag1_7 : _GEN_10; // @[DCache.scala 63:28 DCache.scala 63:28]
  wire [52:0] _GEN_12 = 5'h8 == index_addr ? tag1_8 : _GEN_11; // @[DCache.scala 63:28 DCache.scala 63:28]
  wire [52:0] _GEN_13 = 5'h9 == index_addr ? tag1_9 : _GEN_12; // @[DCache.scala 63:28 DCache.scala 63:28]
  wire [52:0] _GEN_14 = 5'ha == index_addr ? tag1_10 : _GEN_13; // @[DCache.scala 63:28 DCache.scala 63:28]
  wire [52:0] _GEN_15 = 5'hb == index_addr ? tag1_11 : _GEN_14; // @[DCache.scala 63:28 DCache.scala 63:28]
  wire [52:0] _GEN_16 = 5'hc == index_addr ? tag1_12 : _GEN_15; // @[DCache.scala 63:28 DCache.scala 63:28]
  wire [52:0] _GEN_17 = 5'hd == index_addr ? tag1_13 : _GEN_16; // @[DCache.scala 63:28 DCache.scala 63:28]
  wire [52:0] _GEN_18 = 5'he == index_addr ? tag1_14 : _GEN_17; // @[DCache.scala 63:28 DCache.scala 63:28]
  wire [52:0] _GEN_19 = 5'hf == index_addr ? tag1_15 : _GEN_18; // @[DCache.scala 63:28 DCache.scala 63:28]
  wire [52:0] _GEN_20 = 5'h10 == index_addr ? tag1_16 : _GEN_19; // @[DCache.scala 63:28 DCache.scala 63:28]
  wire [52:0] _GEN_21 = 5'h11 == index_addr ? tag1_17 : _GEN_20; // @[DCache.scala 63:28 DCache.scala 63:28]
  wire [52:0] _GEN_22 = 5'h12 == index_addr ? tag1_18 : _GEN_21; // @[DCache.scala 63:28 DCache.scala 63:28]
  wire [52:0] _GEN_23 = 5'h13 == index_addr ? tag1_19 : _GEN_22; // @[DCache.scala 63:28 DCache.scala 63:28]
  wire [52:0] _GEN_24 = 5'h14 == index_addr ? tag1_20 : _GEN_23; // @[DCache.scala 63:28 DCache.scala 63:28]
  wire [52:0] _GEN_25 = 5'h15 == index_addr ? tag1_21 : _GEN_24; // @[DCache.scala 63:28 DCache.scala 63:28]
  wire [52:0] _GEN_26 = 5'h16 == index_addr ? tag1_22 : _GEN_25; // @[DCache.scala 63:28 DCache.scala 63:28]
  wire [52:0] _GEN_27 = 5'h17 == index_addr ? tag1_23 : _GEN_26; // @[DCache.scala 63:28 DCache.scala 63:28]
  wire [52:0] _GEN_28 = 5'h18 == index_addr ? tag1_24 : _GEN_27; // @[DCache.scala 63:28 DCache.scala 63:28]
  wire [52:0] _GEN_29 = 5'h19 == index_addr ? tag1_25 : _GEN_28; // @[DCache.scala 63:28 DCache.scala 63:28]
  wire [52:0] _GEN_30 = 5'h1a == index_addr ? tag1_26 : _GEN_29; // @[DCache.scala 63:28 DCache.scala 63:28]
  wire [52:0] _GEN_31 = 5'h1b == index_addr ? tag1_27 : _GEN_30; // @[DCache.scala 63:28 DCache.scala 63:28]
  wire [52:0] _GEN_32 = 5'h1c == index_addr ? tag1_28 : _GEN_31; // @[DCache.scala 63:28 DCache.scala 63:28]
  wire [52:0] _GEN_33 = 5'h1d == index_addr ? tag1_29 : _GEN_32; // @[DCache.scala 63:28 DCache.scala 63:28]
  wire [52:0] _GEN_34 = 5'h1e == index_addr ? tag1_30 : _GEN_33; // @[DCache.scala 63:28 DCache.scala 63:28]
  wire [52:0] _GEN_35 = 5'h1f == index_addr ? tag1_31 : _GEN_34; // @[DCache.scala 63:28 DCache.scala 63:28]
  wire  _GEN_37 = 5'h1 == index_addr ? v1_1 : v1_0; // @[DCache.scala 63:67 DCache.scala 63:67]
  wire  _GEN_38 = 5'h2 == index_addr ? v1_2 : _GEN_37; // @[DCache.scala 63:67 DCache.scala 63:67]
  wire  _GEN_39 = 5'h3 == index_addr ? v1_3 : _GEN_38; // @[DCache.scala 63:67 DCache.scala 63:67]
  wire  _GEN_40 = 5'h4 == index_addr ? v1_4 : _GEN_39; // @[DCache.scala 63:67 DCache.scala 63:67]
  wire  _GEN_41 = 5'h5 == index_addr ? v1_5 : _GEN_40; // @[DCache.scala 63:67 DCache.scala 63:67]
  wire  _GEN_42 = 5'h6 == index_addr ? v1_6 : _GEN_41; // @[DCache.scala 63:67 DCache.scala 63:67]
  wire  _GEN_43 = 5'h7 == index_addr ? v1_7 : _GEN_42; // @[DCache.scala 63:67 DCache.scala 63:67]
  wire  _GEN_44 = 5'h8 == index_addr ? v1_8 : _GEN_43; // @[DCache.scala 63:67 DCache.scala 63:67]
  wire  _GEN_45 = 5'h9 == index_addr ? v1_9 : _GEN_44; // @[DCache.scala 63:67 DCache.scala 63:67]
  wire  _GEN_46 = 5'ha == index_addr ? v1_10 : _GEN_45; // @[DCache.scala 63:67 DCache.scala 63:67]
  wire  _GEN_47 = 5'hb == index_addr ? v1_11 : _GEN_46; // @[DCache.scala 63:67 DCache.scala 63:67]
  wire  _GEN_48 = 5'hc == index_addr ? v1_12 : _GEN_47; // @[DCache.scala 63:67 DCache.scala 63:67]
  wire  _GEN_49 = 5'hd == index_addr ? v1_13 : _GEN_48; // @[DCache.scala 63:67 DCache.scala 63:67]
  wire  _GEN_50 = 5'he == index_addr ? v1_14 : _GEN_49; // @[DCache.scala 63:67 DCache.scala 63:67]
  wire  _GEN_51 = 5'hf == index_addr ? v1_15 : _GEN_50; // @[DCache.scala 63:67 DCache.scala 63:67]
  wire  _GEN_52 = 5'h10 == index_addr ? v1_16 : _GEN_51; // @[DCache.scala 63:67 DCache.scala 63:67]
  wire  _GEN_53 = 5'h11 == index_addr ? v1_17 : _GEN_52; // @[DCache.scala 63:67 DCache.scala 63:67]
  wire  _GEN_54 = 5'h12 == index_addr ? v1_18 : _GEN_53; // @[DCache.scala 63:67 DCache.scala 63:67]
  wire  _GEN_55 = 5'h13 == index_addr ? v1_19 : _GEN_54; // @[DCache.scala 63:67 DCache.scala 63:67]
  wire  _GEN_56 = 5'h14 == index_addr ? v1_20 : _GEN_55; // @[DCache.scala 63:67 DCache.scala 63:67]
  wire  _GEN_57 = 5'h15 == index_addr ? v1_21 : _GEN_56; // @[DCache.scala 63:67 DCache.scala 63:67]
  wire  _GEN_58 = 5'h16 == index_addr ? v1_22 : _GEN_57; // @[DCache.scala 63:67 DCache.scala 63:67]
  wire  _GEN_59 = 5'h17 == index_addr ? v1_23 : _GEN_58; // @[DCache.scala 63:67 DCache.scala 63:67]
  wire  _GEN_60 = 5'h18 == index_addr ? v1_24 : _GEN_59; // @[DCache.scala 63:67 DCache.scala 63:67]
  wire  _GEN_61 = 5'h19 == index_addr ? v1_25 : _GEN_60; // @[DCache.scala 63:67 DCache.scala 63:67]
  wire  _GEN_62 = 5'h1a == index_addr ? v1_26 : _GEN_61; // @[DCache.scala 63:67 DCache.scala 63:67]
  wire  _GEN_63 = 5'h1b == index_addr ? v1_27 : _GEN_62; // @[DCache.scala 63:67 DCache.scala 63:67]
  wire  _GEN_64 = 5'h1c == index_addr ? v1_28 : _GEN_63; // @[DCache.scala 63:67 DCache.scala 63:67]
  wire  _GEN_65 = 5'h1d == index_addr ? v1_29 : _GEN_64; // @[DCache.scala 63:67 DCache.scala 63:67]
  wire  _GEN_66 = 5'h1e == index_addr ? v1_30 : _GEN_65; // @[DCache.scala 63:67 DCache.scala 63:67]
  wire  _GEN_67 = 5'h1f == index_addr ? v1_31 : _GEN_66; // @[DCache.scala 63:67 DCache.scala 63:67]
  wire  hit1 = tag_addr == _GEN_35 & _GEN_67; // @[DCache.scala 63:49]
  wire [52:0] _GEN_69 = 5'h1 == index_addr ? tag2_1 : tag2_0; // @[DCache.scala 64:28 DCache.scala 64:28]
  wire [52:0] _GEN_70 = 5'h2 == index_addr ? tag2_2 : _GEN_69; // @[DCache.scala 64:28 DCache.scala 64:28]
  wire [52:0] _GEN_71 = 5'h3 == index_addr ? tag2_3 : _GEN_70; // @[DCache.scala 64:28 DCache.scala 64:28]
  wire [52:0] _GEN_72 = 5'h4 == index_addr ? tag2_4 : _GEN_71; // @[DCache.scala 64:28 DCache.scala 64:28]
  wire [52:0] _GEN_73 = 5'h5 == index_addr ? tag2_5 : _GEN_72; // @[DCache.scala 64:28 DCache.scala 64:28]
  wire [52:0] _GEN_74 = 5'h6 == index_addr ? tag2_6 : _GEN_73; // @[DCache.scala 64:28 DCache.scala 64:28]
  wire [52:0] _GEN_75 = 5'h7 == index_addr ? tag2_7 : _GEN_74; // @[DCache.scala 64:28 DCache.scala 64:28]
  wire [52:0] _GEN_76 = 5'h8 == index_addr ? tag2_8 : _GEN_75; // @[DCache.scala 64:28 DCache.scala 64:28]
  wire [52:0] _GEN_77 = 5'h9 == index_addr ? tag2_9 : _GEN_76; // @[DCache.scala 64:28 DCache.scala 64:28]
  wire [52:0] _GEN_78 = 5'ha == index_addr ? tag2_10 : _GEN_77; // @[DCache.scala 64:28 DCache.scala 64:28]
  wire [52:0] _GEN_79 = 5'hb == index_addr ? tag2_11 : _GEN_78; // @[DCache.scala 64:28 DCache.scala 64:28]
  wire [52:0] _GEN_80 = 5'hc == index_addr ? tag2_12 : _GEN_79; // @[DCache.scala 64:28 DCache.scala 64:28]
  wire [52:0] _GEN_81 = 5'hd == index_addr ? tag2_13 : _GEN_80; // @[DCache.scala 64:28 DCache.scala 64:28]
  wire [52:0] _GEN_82 = 5'he == index_addr ? tag2_14 : _GEN_81; // @[DCache.scala 64:28 DCache.scala 64:28]
  wire [52:0] _GEN_83 = 5'hf == index_addr ? tag2_15 : _GEN_82; // @[DCache.scala 64:28 DCache.scala 64:28]
  wire [52:0] _GEN_84 = 5'h10 == index_addr ? tag2_16 : _GEN_83; // @[DCache.scala 64:28 DCache.scala 64:28]
  wire [52:0] _GEN_85 = 5'h11 == index_addr ? tag2_17 : _GEN_84; // @[DCache.scala 64:28 DCache.scala 64:28]
  wire [52:0] _GEN_86 = 5'h12 == index_addr ? tag2_18 : _GEN_85; // @[DCache.scala 64:28 DCache.scala 64:28]
  wire [52:0] _GEN_87 = 5'h13 == index_addr ? tag2_19 : _GEN_86; // @[DCache.scala 64:28 DCache.scala 64:28]
  wire [52:0] _GEN_88 = 5'h14 == index_addr ? tag2_20 : _GEN_87; // @[DCache.scala 64:28 DCache.scala 64:28]
  wire [52:0] _GEN_89 = 5'h15 == index_addr ? tag2_21 : _GEN_88; // @[DCache.scala 64:28 DCache.scala 64:28]
  wire [52:0] _GEN_90 = 5'h16 == index_addr ? tag2_22 : _GEN_89; // @[DCache.scala 64:28 DCache.scala 64:28]
  wire [52:0] _GEN_91 = 5'h17 == index_addr ? tag2_23 : _GEN_90; // @[DCache.scala 64:28 DCache.scala 64:28]
  wire [52:0] _GEN_92 = 5'h18 == index_addr ? tag2_24 : _GEN_91; // @[DCache.scala 64:28 DCache.scala 64:28]
  wire [52:0] _GEN_93 = 5'h19 == index_addr ? tag2_25 : _GEN_92; // @[DCache.scala 64:28 DCache.scala 64:28]
  wire [52:0] _GEN_94 = 5'h1a == index_addr ? tag2_26 : _GEN_93; // @[DCache.scala 64:28 DCache.scala 64:28]
  wire [52:0] _GEN_95 = 5'h1b == index_addr ? tag2_27 : _GEN_94; // @[DCache.scala 64:28 DCache.scala 64:28]
  wire [52:0] _GEN_96 = 5'h1c == index_addr ? tag2_28 : _GEN_95; // @[DCache.scala 64:28 DCache.scala 64:28]
  wire [52:0] _GEN_97 = 5'h1d == index_addr ? tag2_29 : _GEN_96; // @[DCache.scala 64:28 DCache.scala 64:28]
  wire [52:0] _GEN_98 = 5'h1e == index_addr ? tag2_30 : _GEN_97; // @[DCache.scala 64:28 DCache.scala 64:28]
  wire [52:0] _GEN_99 = 5'h1f == index_addr ? tag2_31 : _GEN_98; // @[DCache.scala 64:28 DCache.scala 64:28]
  wire  _GEN_101 = 5'h1 == index_addr ? v2_1 : v2_0; // @[DCache.scala 64:67 DCache.scala 64:67]
  wire  _GEN_102 = 5'h2 == index_addr ? v2_2 : _GEN_101; // @[DCache.scala 64:67 DCache.scala 64:67]
  wire  _GEN_103 = 5'h3 == index_addr ? v2_3 : _GEN_102; // @[DCache.scala 64:67 DCache.scala 64:67]
  wire  _GEN_104 = 5'h4 == index_addr ? v2_4 : _GEN_103; // @[DCache.scala 64:67 DCache.scala 64:67]
  wire  _GEN_105 = 5'h5 == index_addr ? v2_5 : _GEN_104; // @[DCache.scala 64:67 DCache.scala 64:67]
  wire  _GEN_106 = 5'h6 == index_addr ? v2_6 : _GEN_105; // @[DCache.scala 64:67 DCache.scala 64:67]
  wire  _GEN_107 = 5'h7 == index_addr ? v2_7 : _GEN_106; // @[DCache.scala 64:67 DCache.scala 64:67]
  wire  _GEN_108 = 5'h8 == index_addr ? v2_8 : _GEN_107; // @[DCache.scala 64:67 DCache.scala 64:67]
  wire  _GEN_109 = 5'h9 == index_addr ? v2_9 : _GEN_108; // @[DCache.scala 64:67 DCache.scala 64:67]
  wire  _GEN_110 = 5'ha == index_addr ? v2_10 : _GEN_109; // @[DCache.scala 64:67 DCache.scala 64:67]
  wire  _GEN_111 = 5'hb == index_addr ? v2_11 : _GEN_110; // @[DCache.scala 64:67 DCache.scala 64:67]
  wire  _GEN_112 = 5'hc == index_addr ? v2_12 : _GEN_111; // @[DCache.scala 64:67 DCache.scala 64:67]
  wire  _GEN_113 = 5'hd == index_addr ? v2_13 : _GEN_112; // @[DCache.scala 64:67 DCache.scala 64:67]
  wire  _GEN_114 = 5'he == index_addr ? v2_14 : _GEN_113; // @[DCache.scala 64:67 DCache.scala 64:67]
  wire  _GEN_115 = 5'hf == index_addr ? v2_15 : _GEN_114; // @[DCache.scala 64:67 DCache.scala 64:67]
  wire  _GEN_116 = 5'h10 == index_addr ? v2_16 : _GEN_115; // @[DCache.scala 64:67 DCache.scala 64:67]
  wire  _GEN_117 = 5'h11 == index_addr ? v2_17 : _GEN_116; // @[DCache.scala 64:67 DCache.scala 64:67]
  wire  _GEN_118 = 5'h12 == index_addr ? v2_18 : _GEN_117; // @[DCache.scala 64:67 DCache.scala 64:67]
  wire  _GEN_119 = 5'h13 == index_addr ? v2_19 : _GEN_118; // @[DCache.scala 64:67 DCache.scala 64:67]
  wire  _GEN_120 = 5'h14 == index_addr ? v2_20 : _GEN_119; // @[DCache.scala 64:67 DCache.scala 64:67]
  wire  _GEN_121 = 5'h15 == index_addr ? v2_21 : _GEN_120; // @[DCache.scala 64:67 DCache.scala 64:67]
  wire  _GEN_122 = 5'h16 == index_addr ? v2_22 : _GEN_121; // @[DCache.scala 64:67 DCache.scala 64:67]
  wire  _GEN_123 = 5'h17 == index_addr ? v2_23 : _GEN_122; // @[DCache.scala 64:67 DCache.scala 64:67]
  wire  _GEN_124 = 5'h18 == index_addr ? v2_24 : _GEN_123; // @[DCache.scala 64:67 DCache.scala 64:67]
  wire  _GEN_125 = 5'h19 == index_addr ? v2_25 : _GEN_124; // @[DCache.scala 64:67 DCache.scala 64:67]
  wire  _GEN_126 = 5'h1a == index_addr ? v2_26 : _GEN_125; // @[DCache.scala 64:67 DCache.scala 64:67]
  wire  _GEN_127 = 5'h1b == index_addr ? v2_27 : _GEN_126; // @[DCache.scala 64:67 DCache.scala 64:67]
  wire  _GEN_128 = 5'h1c == index_addr ? v2_28 : _GEN_127; // @[DCache.scala 64:67 DCache.scala 64:67]
  wire  _GEN_129 = 5'h1d == index_addr ? v2_29 : _GEN_128; // @[DCache.scala 64:67 DCache.scala 64:67]
  wire  _GEN_130 = 5'h1e == index_addr ? v2_30 : _GEN_129; // @[DCache.scala 64:67 DCache.scala 64:67]
  wire  _GEN_131 = 5'h1f == index_addr ? v2_31 : _GEN_130; // @[DCache.scala 64:67 DCache.scala 64:67]
  wire  hit2 = tag_addr == _GEN_99 & _GEN_131; // @[DCache.scala 64:49]
  wire [8:0] _rdata1_T = {offset_addr, 3'h0}; // @[DCache.scala 65:55]
  wire [511:0] _GEN_133 = 5'h1 == index_addr ? block1_1 : block1_0; // @[DCache.scala 65:39 DCache.scala 65:39]
  wire [511:0] _GEN_134 = 5'h2 == index_addr ? block1_2 : _GEN_133; // @[DCache.scala 65:39 DCache.scala 65:39]
  wire [511:0] _GEN_135 = 5'h3 == index_addr ? block1_3 : _GEN_134; // @[DCache.scala 65:39 DCache.scala 65:39]
  wire [511:0] _GEN_136 = 5'h4 == index_addr ? block1_4 : _GEN_135; // @[DCache.scala 65:39 DCache.scala 65:39]
  wire [511:0] _GEN_137 = 5'h5 == index_addr ? block1_5 : _GEN_136; // @[DCache.scala 65:39 DCache.scala 65:39]
  wire [511:0] _GEN_138 = 5'h6 == index_addr ? block1_6 : _GEN_137; // @[DCache.scala 65:39 DCache.scala 65:39]
  wire [511:0] _GEN_139 = 5'h7 == index_addr ? block1_7 : _GEN_138; // @[DCache.scala 65:39 DCache.scala 65:39]
  wire [511:0] _GEN_140 = 5'h8 == index_addr ? block1_8 : _GEN_139; // @[DCache.scala 65:39 DCache.scala 65:39]
  wire [511:0] _GEN_141 = 5'h9 == index_addr ? block1_9 : _GEN_140; // @[DCache.scala 65:39 DCache.scala 65:39]
  wire [511:0] _GEN_142 = 5'ha == index_addr ? block1_10 : _GEN_141; // @[DCache.scala 65:39 DCache.scala 65:39]
  wire [511:0] _GEN_143 = 5'hb == index_addr ? block1_11 : _GEN_142; // @[DCache.scala 65:39 DCache.scala 65:39]
  wire [511:0] _GEN_144 = 5'hc == index_addr ? block1_12 : _GEN_143; // @[DCache.scala 65:39 DCache.scala 65:39]
  wire [511:0] _GEN_145 = 5'hd == index_addr ? block1_13 : _GEN_144; // @[DCache.scala 65:39 DCache.scala 65:39]
  wire [511:0] _GEN_146 = 5'he == index_addr ? block1_14 : _GEN_145; // @[DCache.scala 65:39 DCache.scala 65:39]
  wire [511:0] _GEN_147 = 5'hf == index_addr ? block1_15 : _GEN_146; // @[DCache.scala 65:39 DCache.scala 65:39]
  wire [511:0] _GEN_148 = 5'h10 == index_addr ? block1_16 : _GEN_147; // @[DCache.scala 65:39 DCache.scala 65:39]
  wire [511:0] _GEN_149 = 5'h11 == index_addr ? block1_17 : _GEN_148; // @[DCache.scala 65:39 DCache.scala 65:39]
  wire [511:0] _GEN_150 = 5'h12 == index_addr ? block1_18 : _GEN_149; // @[DCache.scala 65:39 DCache.scala 65:39]
  wire [511:0] _GEN_151 = 5'h13 == index_addr ? block1_19 : _GEN_150; // @[DCache.scala 65:39 DCache.scala 65:39]
  wire [511:0] _GEN_152 = 5'h14 == index_addr ? block1_20 : _GEN_151; // @[DCache.scala 65:39 DCache.scala 65:39]
  wire [511:0] _GEN_153 = 5'h15 == index_addr ? block1_21 : _GEN_152; // @[DCache.scala 65:39 DCache.scala 65:39]
  wire [511:0] _GEN_154 = 5'h16 == index_addr ? block1_22 : _GEN_153; // @[DCache.scala 65:39 DCache.scala 65:39]
  wire [511:0] _GEN_155 = 5'h17 == index_addr ? block1_23 : _GEN_154; // @[DCache.scala 65:39 DCache.scala 65:39]
  wire [511:0] _GEN_156 = 5'h18 == index_addr ? block1_24 : _GEN_155; // @[DCache.scala 65:39 DCache.scala 65:39]
  wire [511:0] _GEN_157 = 5'h19 == index_addr ? block1_25 : _GEN_156; // @[DCache.scala 65:39 DCache.scala 65:39]
  wire [511:0] _GEN_158 = 5'h1a == index_addr ? block1_26 : _GEN_157; // @[DCache.scala 65:39 DCache.scala 65:39]
  wire [511:0] _GEN_159 = 5'h1b == index_addr ? block1_27 : _GEN_158; // @[DCache.scala 65:39 DCache.scala 65:39]
  wire [511:0] _GEN_160 = 5'h1c == index_addr ? block1_28 : _GEN_159; // @[DCache.scala 65:39 DCache.scala 65:39]
  wire [511:0] _GEN_161 = 5'h1d == index_addr ? block1_29 : _GEN_160; // @[DCache.scala 65:39 DCache.scala 65:39]
  wire [511:0] _GEN_162 = 5'h1e == index_addr ? block1_30 : _GEN_161; // @[DCache.scala 65:39 DCache.scala 65:39]
  wire [511:0] _GEN_163 = 5'h1f == index_addr ? block1_31 : _GEN_162; // @[DCache.scala 65:39 DCache.scala 65:39]
  wire [511:0] _rdata1_T_1 = _GEN_163 >> _rdata1_T; // @[DCache.scala 65:39]
  wire [63:0] rdata1 = _rdata1_T_1[63:0]; // @[DCache.scala 65:61]
  wire [511:0] _GEN_165 = 5'h1 == index_addr ? block2_1 : block2_0; // @[DCache.scala 66:39 DCache.scala 66:39]
  wire [511:0] _GEN_166 = 5'h2 == index_addr ? block2_2 : _GEN_165; // @[DCache.scala 66:39 DCache.scala 66:39]
  wire [511:0] _GEN_167 = 5'h3 == index_addr ? block2_3 : _GEN_166; // @[DCache.scala 66:39 DCache.scala 66:39]
  wire [511:0] _GEN_168 = 5'h4 == index_addr ? block2_4 : _GEN_167; // @[DCache.scala 66:39 DCache.scala 66:39]
  wire [511:0] _GEN_169 = 5'h5 == index_addr ? block2_5 : _GEN_168; // @[DCache.scala 66:39 DCache.scala 66:39]
  wire [511:0] _GEN_170 = 5'h6 == index_addr ? block2_6 : _GEN_169; // @[DCache.scala 66:39 DCache.scala 66:39]
  wire [511:0] _GEN_171 = 5'h7 == index_addr ? block2_7 : _GEN_170; // @[DCache.scala 66:39 DCache.scala 66:39]
  wire [511:0] _GEN_172 = 5'h8 == index_addr ? block2_8 : _GEN_171; // @[DCache.scala 66:39 DCache.scala 66:39]
  wire [511:0] _GEN_173 = 5'h9 == index_addr ? block2_9 : _GEN_172; // @[DCache.scala 66:39 DCache.scala 66:39]
  wire [511:0] _GEN_174 = 5'ha == index_addr ? block2_10 : _GEN_173; // @[DCache.scala 66:39 DCache.scala 66:39]
  wire [511:0] _GEN_175 = 5'hb == index_addr ? block2_11 : _GEN_174; // @[DCache.scala 66:39 DCache.scala 66:39]
  wire [511:0] _GEN_176 = 5'hc == index_addr ? block2_12 : _GEN_175; // @[DCache.scala 66:39 DCache.scala 66:39]
  wire [511:0] _GEN_177 = 5'hd == index_addr ? block2_13 : _GEN_176; // @[DCache.scala 66:39 DCache.scala 66:39]
  wire [511:0] _GEN_178 = 5'he == index_addr ? block2_14 : _GEN_177; // @[DCache.scala 66:39 DCache.scala 66:39]
  wire [511:0] _GEN_179 = 5'hf == index_addr ? block2_15 : _GEN_178; // @[DCache.scala 66:39 DCache.scala 66:39]
  wire [511:0] _GEN_180 = 5'h10 == index_addr ? block2_16 : _GEN_179; // @[DCache.scala 66:39 DCache.scala 66:39]
  wire [511:0] _GEN_181 = 5'h11 == index_addr ? block2_17 : _GEN_180; // @[DCache.scala 66:39 DCache.scala 66:39]
  wire [511:0] _GEN_182 = 5'h12 == index_addr ? block2_18 : _GEN_181; // @[DCache.scala 66:39 DCache.scala 66:39]
  wire [511:0] _GEN_183 = 5'h13 == index_addr ? block2_19 : _GEN_182; // @[DCache.scala 66:39 DCache.scala 66:39]
  wire [511:0] _GEN_184 = 5'h14 == index_addr ? block2_20 : _GEN_183; // @[DCache.scala 66:39 DCache.scala 66:39]
  wire [511:0] _GEN_185 = 5'h15 == index_addr ? block2_21 : _GEN_184; // @[DCache.scala 66:39 DCache.scala 66:39]
  wire [511:0] _GEN_186 = 5'h16 == index_addr ? block2_22 : _GEN_185; // @[DCache.scala 66:39 DCache.scala 66:39]
  wire [511:0] _GEN_187 = 5'h17 == index_addr ? block2_23 : _GEN_186; // @[DCache.scala 66:39 DCache.scala 66:39]
  wire [511:0] _GEN_188 = 5'h18 == index_addr ? block2_24 : _GEN_187; // @[DCache.scala 66:39 DCache.scala 66:39]
  wire [511:0] _GEN_189 = 5'h19 == index_addr ? block2_25 : _GEN_188; // @[DCache.scala 66:39 DCache.scala 66:39]
  wire [511:0] _GEN_190 = 5'h1a == index_addr ? block2_26 : _GEN_189; // @[DCache.scala 66:39 DCache.scala 66:39]
  wire [511:0] _GEN_191 = 5'h1b == index_addr ? block2_27 : _GEN_190; // @[DCache.scala 66:39 DCache.scala 66:39]
  wire [511:0] _GEN_192 = 5'h1c == index_addr ? block2_28 : _GEN_191; // @[DCache.scala 66:39 DCache.scala 66:39]
  wire [511:0] _GEN_193 = 5'h1d == index_addr ? block2_29 : _GEN_192; // @[DCache.scala 66:39 DCache.scala 66:39]
  wire [511:0] _GEN_194 = 5'h1e == index_addr ? block2_30 : _GEN_193; // @[DCache.scala 66:39 DCache.scala 66:39]
  wire [511:0] _GEN_195 = 5'h1f == index_addr ? block2_31 : _GEN_194; // @[DCache.scala 66:39 DCache.scala 66:39]
  wire [511:0] _rdata2_T_1 = _GEN_195 >> _rdata1_T; // @[DCache.scala 66:39]
  wire [63:0] rdata2 = _rdata2_T_1[63:0]; // @[DCache.scala 66:61]
  reg [2:0] state; // @[DCache.scala 69:24]
  wire  hit = hit1 | hit2; // @[DCache.scala 71:28]
  wire [63:0] _rdata_T = hit1 ? rdata1 : 64'h0; // @[DCache.scala 72:44]
  reg  not_en_yet; // @[DCache.scala 74:30]
  wire  _not_en_yet_T = io_dmem_en ? 1'h0 : not_en_yet; // @[DCache.scala 75:27]
  wire  _age1_T = hit1 ^ hit2; // @[DCache.scala 81:35]
  wire  _GEN_197 = 5'h1 == index_addr ? age1_1 : age1_0; // @[DCache.scala 81:28 DCache.scala 81:28]
  wire  _GEN_198 = 5'h2 == index_addr ? age1_2 : _GEN_197; // @[DCache.scala 81:28 DCache.scala 81:28]
  wire  _GEN_199 = 5'h3 == index_addr ? age1_3 : _GEN_198; // @[DCache.scala 81:28 DCache.scala 81:28]
  wire  _GEN_200 = 5'h4 == index_addr ? age1_4 : _GEN_199; // @[DCache.scala 81:28 DCache.scala 81:28]
  wire  _GEN_201 = 5'h5 == index_addr ? age1_5 : _GEN_200; // @[DCache.scala 81:28 DCache.scala 81:28]
  wire  _GEN_202 = 5'h6 == index_addr ? age1_6 : _GEN_201; // @[DCache.scala 81:28 DCache.scala 81:28]
  wire  _GEN_203 = 5'h7 == index_addr ? age1_7 : _GEN_202; // @[DCache.scala 81:28 DCache.scala 81:28]
  wire  _GEN_204 = 5'h8 == index_addr ? age1_8 : _GEN_203; // @[DCache.scala 81:28 DCache.scala 81:28]
  wire  _GEN_205 = 5'h9 == index_addr ? age1_9 : _GEN_204; // @[DCache.scala 81:28 DCache.scala 81:28]
  wire  _GEN_206 = 5'ha == index_addr ? age1_10 : _GEN_205; // @[DCache.scala 81:28 DCache.scala 81:28]
  wire  _GEN_207 = 5'hb == index_addr ? age1_11 : _GEN_206; // @[DCache.scala 81:28 DCache.scala 81:28]
  wire  _GEN_208 = 5'hc == index_addr ? age1_12 : _GEN_207; // @[DCache.scala 81:28 DCache.scala 81:28]
  wire  _GEN_209 = 5'hd == index_addr ? age1_13 : _GEN_208; // @[DCache.scala 81:28 DCache.scala 81:28]
  wire  _GEN_210 = 5'he == index_addr ? age1_14 : _GEN_209; // @[DCache.scala 81:28 DCache.scala 81:28]
  wire  _GEN_211 = 5'hf == index_addr ? age1_15 : _GEN_210; // @[DCache.scala 81:28 DCache.scala 81:28]
  wire  _GEN_212 = 5'h10 == index_addr ? age1_16 : _GEN_211; // @[DCache.scala 81:28 DCache.scala 81:28]
  wire  _GEN_213 = 5'h11 == index_addr ? age1_17 : _GEN_212; // @[DCache.scala 81:28 DCache.scala 81:28]
  wire  _GEN_214 = 5'h12 == index_addr ? age1_18 : _GEN_213; // @[DCache.scala 81:28 DCache.scala 81:28]
  wire  _GEN_215 = 5'h13 == index_addr ? age1_19 : _GEN_214; // @[DCache.scala 81:28 DCache.scala 81:28]
  wire  _GEN_216 = 5'h14 == index_addr ? age1_20 : _GEN_215; // @[DCache.scala 81:28 DCache.scala 81:28]
  wire  _GEN_217 = 5'h15 == index_addr ? age1_21 : _GEN_216; // @[DCache.scala 81:28 DCache.scala 81:28]
  wire  _GEN_218 = 5'h16 == index_addr ? age1_22 : _GEN_217; // @[DCache.scala 81:28 DCache.scala 81:28]
  wire  _GEN_219 = 5'h17 == index_addr ? age1_23 : _GEN_218; // @[DCache.scala 81:28 DCache.scala 81:28]
  wire  _GEN_220 = 5'h18 == index_addr ? age1_24 : _GEN_219; // @[DCache.scala 81:28 DCache.scala 81:28]
  wire  _GEN_221 = 5'h19 == index_addr ? age1_25 : _GEN_220; // @[DCache.scala 81:28 DCache.scala 81:28]
  wire  _GEN_222 = 5'h1a == index_addr ? age1_26 : _GEN_221; // @[DCache.scala 81:28 DCache.scala 81:28]
  wire  _GEN_223 = 5'h1b == index_addr ? age1_27 : _GEN_222; // @[DCache.scala 81:28 DCache.scala 81:28]
  wire  _GEN_224 = 5'h1c == index_addr ? age1_28 : _GEN_223; // @[DCache.scala 81:28 DCache.scala 81:28]
  wire  _GEN_225 = 5'h1d == index_addr ? age1_29 : _GEN_224; // @[DCache.scala 81:28 DCache.scala 81:28]
  wire  _GEN_226 = 5'h1e == index_addr ? age1_30 : _GEN_225; // @[DCache.scala 81:28 DCache.scala 81:28]
  wire  _GEN_227 = 5'h1f == index_addr ? age1_31 : _GEN_226; // @[DCache.scala 81:28 DCache.scala 81:28]
  wire  _GEN_261 = 5'h1 == index_addr ? age2_1 : age2_0; // @[DCache.scala 82:28 DCache.scala 82:28]
  wire  _GEN_262 = 5'h2 == index_addr ? age2_2 : _GEN_261; // @[DCache.scala 82:28 DCache.scala 82:28]
  wire  _GEN_263 = 5'h3 == index_addr ? age2_3 : _GEN_262; // @[DCache.scala 82:28 DCache.scala 82:28]
  wire  _GEN_264 = 5'h4 == index_addr ? age2_4 : _GEN_263; // @[DCache.scala 82:28 DCache.scala 82:28]
  wire  _GEN_265 = 5'h5 == index_addr ? age2_5 : _GEN_264; // @[DCache.scala 82:28 DCache.scala 82:28]
  wire  _GEN_266 = 5'h6 == index_addr ? age2_6 : _GEN_265; // @[DCache.scala 82:28 DCache.scala 82:28]
  wire  _GEN_267 = 5'h7 == index_addr ? age2_7 : _GEN_266; // @[DCache.scala 82:28 DCache.scala 82:28]
  wire  _GEN_268 = 5'h8 == index_addr ? age2_8 : _GEN_267; // @[DCache.scala 82:28 DCache.scala 82:28]
  wire  _GEN_269 = 5'h9 == index_addr ? age2_9 : _GEN_268; // @[DCache.scala 82:28 DCache.scala 82:28]
  wire  _GEN_270 = 5'ha == index_addr ? age2_10 : _GEN_269; // @[DCache.scala 82:28 DCache.scala 82:28]
  wire  _GEN_271 = 5'hb == index_addr ? age2_11 : _GEN_270; // @[DCache.scala 82:28 DCache.scala 82:28]
  wire  _GEN_272 = 5'hc == index_addr ? age2_12 : _GEN_271; // @[DCache.scala 82:28 DCache.scala 82:28]
  wire  _GEN_273 = 5'hd == index_addr ? age2_13 : _GEN_272; // @[DCache.scala 82:28 DCache.scala 82:28]
  wire  _GEN_274 = 5'he == index_addr ? age2_14 : _GEN_273; // @[DCache.scala 82:28 DCache.scala 82:28]
  wire  _GEN_275 = 5'hf == index_addr ? age2_15 : _GEN_274; // @[DCache.scala 82:28 DCache.scala 82:28]
  wire  _GEN_276 = 5'h10 == index_addr ? age2_16 : _GEN_275; // @[DCache.scala 82:28 DCache.scala 82:28]
  wire  _GEN_277 = 5'h11 == index_addr ? age2_17 : _GEN_276; // @[DCache.scala 82:28 DCache.scala 82:28]
  wire  _GEN_278 = 5'h12 == index_addr ? age2_18 : _GEN_277; // @[DCache.scala 82:28 DCache.scala 82:28]
  wire  _GEN_279 = 5'h13 == index_addr ? age2_19 : _GEN_278; // @[DCache.scala 82:28 DCache.scala 82:28]
  wire  _GEN_280 = 5'h14 == index_addr ? age2_20 : _GEN_279; // @[DCache.scala 82:28 DCache.scala 82:28]
  wire  _GEN_281 = 5'h15 == index_addr ? age2_21 : _GEN_280; // @[DCache.scala 82:28 DCache.scala 82:28]
  wire  _GEN_282 = 5'h16 == index_addr ? age2_22 : _GEN_281; // @[DCache.scala 82:28 DCache.scala 82:28]
  wire  _GEN_283 = 5'h17 == index_addr ? age2_23 : _GEN_282; // @[DCache.scala 82:28 DCache.scala 82:28]
  wire  _GEN_284 = 5'h18 == index_addr ? age2_24 : _GEN_283; // @[DCache.scala 82:28 DCache.scala 82:28]
  wire  _GEN_285 = 5'h19 == index_addr ? age2_25 : _GEN_284; // @[DCache.scala 82:28 DCache.scala 82:28]
  wire  _GEN_286 = 5'h1a == index_addr ? age2_26 : _GEN_285; // @[DCache.scala 82:28 DCache.scala 82:28]
  wire  _GEN_287 = 5'h1b == index_addr ? age2_27 : _GEN_286; // @[DCache.scala 82:28 DCache.scala 82:28]
  wire  _GEN_288 = 5'h1c == index_addr ? age2_28 : _GEN_287; // @[DCache.scala 82:28 DCache.scala 82:28]
  wire  _GEN_289 = 5'h1d == index_addr ? age2_29 : _GEN_288; // @[DCache.scala 82:28 DCache.scala 82:28]
  wire  _GEN_290 = 5'h1e == index_addr ? age2_30 : _GEN_289; // @[DCache.scala 82:28 DCache.scala 82:28]
  wire  _GEN_291 = 5'h1f == index_addr ? age2_31 : _GEN_290; // @[DCache.scala 82:28 DCache.scala 82:28]
  wire [1:0] age = {_GEN_291,_GEN_227}; // @[Cat.scala 30:58]
  wire  updateway2 = age == 2'h1; // @[DCache.scala 86:27]
  wire  updateway1 = ~updateway2; // @[DCache.scala 87:23]
  wire  miss = ~hit; // @[DCache.scala 88:23]
  wire  _GEN_325 = 5'h1 == index_addr ? d1_1 : d1_0; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_326 = 5'h2 == index_addr ? d1_2 : _GEN_325; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_327 = 5'h3 == index_addr ? d1_3 : _GEN_326; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_328 = 5'h4 == index_addr ? d1_4 : _GEN_327; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_329 = 5'h5 == index_addr ? d1_5 : _GEN_328; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_330 = 5'h6 == index_addr ? d1_6 : _GEN_329; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_331 = 5'h7 == index_addr ? d1_7 : _GEN_330; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_332 = 5'h8 == index_addr ? d1_8 : _GEN_331; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_333 = 5'h9 == index_addr ? d1_9 : _GEN_332; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_334 = 5'ha == index_addr ? d1_10 : _GEN_333; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_335 = 5'hb == index_addr ? d1_11 : _GEN_334; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_336 = 5'hc == index_addr ? d1_12 : _GEN_335; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_337 = 5'hd == index_addr ? d1_13 : _GEN_336; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_338 = 5'he == index_addr ? d1_14 : _GEN_337; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_339 = 5'hf == index_addr ? d1_15 : _GEN_338; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_340 = 5'h10 == index_addr ? d1_16 : _GEN_339; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_341 = 5'h11 == index_addr ? d1_17 : _GEN_340; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_342 = 5'h12 == index_addr ? d1_18 : _GEN_341; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_343 = 5'h13 == index_addr ? d1_19 : _GEN_342; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_344 = 5'h14 == index_addr ? d1_20 : _GEN_343; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_345 = 5'h15 == index_addr ? d1_21 : _GEN_344; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_346 = 5'h16 == index_addr ? d1_22 : _GEN_345; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_347 = 5'h17 == index_addr ? d1_23 : _GEN_346; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_348 = 5'h18 == index_addr ? d1_24 : _GEN_347; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_349 = 5'h19 == index_addr ? d1_25 : _GEN_348; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_350 = 5'h1a == index_addr ? d1_26 : _GEN_349; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_351 = 5'h1b == index_addr ? d1_27 : _GEN_350; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_352 = 5'h1c == index_addr ? d1_28 : _GEN_351; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_353 = 5'h1d == index_addr ? d1_29 : _GEN_352; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_354 = 5'h1e == index_addr ? d1_30 : _GEN_353; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_355 = 5'h1f == index_addr ? d1_31 : _GEN_354; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_357 = 5'h1 == index_addr ? d2_1 : d2_0; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_358 = 5'h2 == index_addr ? d2_2 : _GEN_357; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_359 = 5'h3 == index_addr ? d2_3 : _GEN_358; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_360 = 5'h4 == index_addr ? d2_4 : _GEN_359; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_361 = 5'h5 == index_addr ? d2_5 : _GEN_360; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_362 = 5'h6 == index_addr ? d2_6 : _GEN_361; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_363 = 5'h7 == index_addr ? d2_7 : _GEN_362; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_364 = 5'h8 == index_addr ? d2_8 : _GEN_363; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_365 = 5'h9 == index_addr ? d2_9 : _GEN_364; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_366 = 5'ha == index_addr ? d2_10 : _GEN_365; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_367 = 5'hb == index_addr ? d2_11 : _GEN_366; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_368 = 5'hc == index_addr ? d2_12 : _GEN_367; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_369 = 5'hd == index_addr ? d2_13 : _GEN_368; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_370 = 5'he == index_addr ? d2_14 : _GEN_369; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_371 = 5'hf == index_addr ? d2_15 : _GEN_370; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_372 = 5'h10 == index_addr ? d2_16 : _GEN_371; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_373 = 5'h11 == index_addr ? d2_17 : _GEN_372; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_374 = 5'h12 == index_addr ? d2_18 : _GEN_373; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_375 = 5'h13 == index_addr ? d2_19 : _GEN_374; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_376 = 5'h14 == index_addr ? d2_20 : _GEN_375; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_377 = 5'h15 == index_addr ? d2_21 : _GEN_376; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_378 = 5'h16 == index_addr ? d2_22 : _GEN_377; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_379 = 5'h17 == index_addr ? d2_23 : _GEN_378; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_380 = 5'h18 == index_addr ? d2_24 : _GEN_379; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_381 = 5'h19 == index_addr ? d2_25 : _GEN_380; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_382 = 5'h1a == index_addr ? d2_26 : _GEN_381; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_383 = 5'h1b == index_addr ? d2_27 : _GEN_382; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_384 = 5'h1c == index_addr ? d2_28 : _GEN_383; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_385 = 5'h1d == index_addr ? d2_29 : _GEN_384; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_386 = 5'h1e == index_addr ? d2_30 : _GEN_385; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  _GEN_387 = 5'h1f == index_addr ? d2_31 : _GEN_386; // @[DCache.scala 89:26 DCache.scala 89:26]
  wire  dirty = updateway1 ? _GEN_355 : _GEN_387; // @[DCache.scala 89:26]
  reg [4:0] fence_cnt; // @[DCache.scala 91:28]
  wire  _T = 3'h0 == state; // @[Conditional.scala 37:30]
  wire [2:0] _state_T = dirty ? 3'h1 : 3'h2; // @[DCache.scala 95:56]
  wire  _T_3 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_4 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_391 = io_axi_rvalid ? 3'h0 : state; // @[DCache.scala 101:33 DCache.scala 101:40 DCache.scala 69:24]
  wire  _T_5 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _GEN_393 = 5'h1 == fence_cnt ? d1_1 : d1_0; // @[DCache.scala 104:32 DCache.scala 104:32]
  wire  _GEN_394 = 5'h2 == fence_cnt ? d1_2 : _GEN_393; // @[DCache.scala 104:32 DCache.scala 104:32]
  wire  _GEN_395 = 5'h3 == fence_cnt ? d1_3 : _GEN_394; // @[DCache.scala 104:32 DCache.scala 104:32]
  wire  _GEN_396 = 5'h4 == fence_cnt ? d1_4 : _GEN_395; // @[DCache.scala 104:32 DCache.scala 104:32]
  wire  _GEN_397 = 5'h5 == fence_cnt ? d1_5 : _GEN_396; // @[DCache.scala 104:32 DCache.scala 104:32]
  wire  _GEN_398 = 5'h6 == fence_cnt ? d1_6 : _GEN_397; // @[DCache.scala 104:32 DCache.scala 104:32]
  wire  _GEN_399 = 5'h7 == fence_cnt ? d1_7 : _GEN_398; // @[DCache.scala 104:32 DCache.scala 104:32]
  wire  _GEN_400 = 5'h8 == fence_cnt ? d1_8 : _GEN_399; // @[DCache.scala 104:32 DCache.scala 104:32]
  wire  _GEN_401 = 5'h9 == fence_cnt ? d1_9 : _GEN_400; // @[DCache.scala 104:32 DCache.scala 104:32]
  wire  _GEN_402 = 5'ha == fence_cnt ? d1_10 : _GEN_401; // @[DCache.scala 104:32 DCache.scala 104:32]
  wire  _GEN_403 = 5'hb == fence_cnt ? d1_11 : _GEN_402; // @[DCache.scala 104:32 DCache.scala 104:32]
  wire  _GEN_404 = 5'hc == fence_cnt ? d1_12 : _GEN_403; // @[DCache.scala 104:32 DCache.scala 104:32]
  wire  _GEN_405 = 5'hd == fence_cnt ? d1_13 : _GEN_404; // @[DCache.scala 104:32 DCache.scala 104:32]
  wire  _GEN_406 = 5'he == fence_cnt ? d1_14 : _GEN_405; // @[DCache.scala 104:32 DCache.scala 104:32]
  wire  _GEN_407 = 5'hf == fence_cnt ? d1_15 : _GEN_406; // @[DCache.scala 104:32 DCache.scala 104:32]
  wire  _GEN_408 = 5'h10 == fence_cnt ? d1_16 : _GEN_407; // @[DCache.scala 104:32 DCache.scala 104:32]
  wire  _GEN_409 = 5'h11 == fence_cnt ? d1_17 : _GEN_408; // @[DCache.scala 104:32 DCache.scala 104:32]
  wire  _GEN_410 = 5'h12 == fence_cnt ? d1_18 : _GEN_409; // @[DCache.scala 104:32 DCache.scala 104:32]
  wire  _GEN_411 = 5'h13 == fence_cnt ? d1_19 : _GEN_410; // @[DCache.scala 104:32 DCache.scala 104:32]
  wire  _GEN_412 = 5'h14 == fence_cnt ? d1_20 : _GEN_411; // @[DCache.scala 104:32 DCache.scala 104:32]
  wire  _GEN_413 = 5'h15 == fence_cnt ? d1_21 : _GEN_412; // @[DCache.scala 104:32 DCache.scala 104:32]
  wire  _GEN_414 = 5'h16 == fence_cnt ? d1_22 : _GEN_413; // @[DCache.scala 104:32 DCache.scala 104:32]
  wire  _GEN_415 = 5'h17 == fence_cnt ? d1_23 : _GEN_414; // @[DCache.scala 104:32 DCache.scala 104:32]
  wire  _GEN_416 = 5'h18 == fence_cnt ? d1_24 : _GEN_415; // @[DCache.scala 104:32 DCache.scala 104:32]
  wire  _GEN_417 = 5'h19 == fence_cnt ? d1_25 : _GEN_416; // @[DCache.scala 104:32 DCache.scala 104:32]
  wire  _GEN_418 = 5'h1a == fence_cnt ? d1_26 : _GEN_417; // @[DCache.scala 104:32 DCache.scala 104:32]
  wire  _GEN_419 = 5'h1b == fence_cnt ? d1_27 : _GEN_418; // @[DCache.scala 104:32 DCache.scala 104:32]
  wire  _GEN_420 = 5'h1c == fence_cnt ? d1_28 : _GEN_419; // @[DCache.scala 104:32 DCache.scala 104:32]
  wire  _GEN_421 = 5'h1d == fence_cnt ? d1_29 : _GEN_420; // @[DCache.scala 104:32 DCache.scala 104:32]
  wire  _GEN_422 = 5'h1e == fence_cnt ? d1_30 : _GEN_421; // @[DCache.scala 104:32 DCache.scala 104:32]
  wire  _GEN_423 = 5'h1f == fence_cnt ? d1_31 : _GEN_422; // @[DCache.scala 104:32 DCache.scala 104:32]
  wire [2:0] _GEN_424 = ~_GEN_423 | _GEN_423 & io_axi_wdone ? 3'h4 : state; // @[DCache.scala 104:91 DCache.scala 104:98 DCache.scala 69:24]
  wire  _T_10 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_11 = fence_cnt == 5'h1f; // @[DCache.scala 107:28]
  wire [2:0] _GEN_425 = fence_cnt == 5'h1f ? 3'h5 : 3'h3; // @[DCache.scala 107:54 DCache.scala 107:61 DCache.scala 108:31]
  wire  _T_12 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_427 = 5'h1 == fence_cnt ? d2_1 : d2_0; // @[DCache.scala 111:32 DCache.scala 111:32]
  wire  _GEN_428 = 5'h2 == fence_cnt ? d2_2 : _GEN_427; // @[DCache.scala 111:32 DCache.scala 111:32]
  wire  _GEN_429 = 5'h3 == fence_cnt ? d2_3 : _GEN_428; // @[DCache.scala 111:32 DCache.scala 111:32]
  wire  _GEN_430 = 5'h4 == fence_cnt ? d2_4 : _GEN_429; // @[DCache.scala 111:32 DCache.scala 111:32]
  wire  _GEN_431 = 5'h5 == fence_cnt ? d2_5 : _GEN_430; // @[DCache.scala 111:32 DCache.scala 111:32]
  wire  _GEN_432 = 5'h6 == fence_cnt ? d2_6 : _GEN_431; // @[DCache.scala 111:32 DCache.scala 111:32]
  wire  _GEN_433 = 5'h7 == fence_cnt ? d2_7 : _GEN_432; // @[DCache.scala 111:32 DCache.scala 111:32]
  wire  _GEN_434 = 5'h8 == fence_cnt ? d2_8 : _GEN_433; // @[DCache.scala 111:32 DCache.scala 111:32]
  wire  _GEN_435 = 5'h9 == fence_cnt ? d2_9 : _GEN_434; // @[DCache.scala 111:32 DCache.scala 111:32]
  wire  _GEN_436 = 5'ha == fence_cnt ? d2_10 : _GEN_435; // @[DCache.scala 111:32 DCache.scala 111:32]
  wire  _GEN_437 = 5'hb == fence_cnt ? d2_11 : _GEN_436; // @[DCache.scala 111:32 DCache.scala 111:32]
  wire  _GEN_438 = 5'hc == fence_cnt ? d2_12 : _GEN_437; // @[DCache.scala 111:32 DCache.scala 111:32]
  wire  _GEN_439 = 5'hd == fence_cnt ? d2_13 : _GEN_438; // @[DCache.scala 111:32 DCache.scala 111:32]
  wire  _GEN_440 = 5'he == fence_cnt ? d2_14 : _GEN_439; // @[DCache.scala 111:32 DCache.scala 111:32]
  wire  _GEN_441 = 5'hf == fence_cnt ? d2_15 : _GEN_440; // @[DCache.scala 111:32 DCache.scala 111:32]
  wire  _GEN_442 = 5'h10 == fence_cnt ? d2_16 : _GEN_441; // @[DCache.scala 111:32 DCache.scala 111:32]
  wire  _GEN_443 = 5'h11 == fence_cnt ? d2_17 : _GEN_442; // @[DCache.scala 111:32 DCache.scala 111:32]
  wire  _GEN_444 = 5'h12 == fence_cnt ? d2_18 : _GEN_443; // @[DCache.scala 111:32 DCache.scala 111:32]
  wire  _GEN_445 = 5'h13 == fence_cnt ? d2_19 : _GEN_444; // @[DCache.scala 111:32 DCache.scala 111:32]
  wire  _GEN_446 = 5'h14 == fence_cnt ? d2_20 : _GEN_445; // @[DCache.scala 111:32 DCache.scala 111:32]
  wire  _GEN_447 = 5'h15 == fence_cnt ? d2_21 : _GEN_446; // @[DCache.scala 111:32 DCache.scala 111:32]
  wire  _GEN_448 = 5'h16 == fence_cnt ? d2_22 : _GEN_447; // @[DCache.scala 111:32 DCache.scala 111:32]
  wire  _GEN_449 = 5'h17 == fence_cnt ? d2_23 : _GEN_448; // @[DCache.scala 111:32 DCache.scala 111:32]
  wire  _GEN_450 = 5'h18 == fence_cnt ? d2_24 : _GEN_449; // @[DCache.scala 111:32 DCache.scala 111:32]
  wire  _GEN_451 = 5'h19 == fence_cnt ? d2_25 : _GEN_450; // @[DCache.scala 111:32 DCache.scala 111:32]
  wire  _GEN_452 = 5'h1a == fence_cnt ? d2_26 : _GEN_451; // @[DCache.scala 111:32 DCache.scala 111:32]
  wire  _GEN_453 = 5'h1b == fence_cnt ? d2_27 : _GEN_452; // @[DCache.scala 111:32 DCache.scala 111:32]
  wire  _GEN_454 = 5'h1c == fence_cnt ? d2_28 : _GEN_453; // @[DCache.scala 111:32 DCache.scala 111:32]
  wire  _GEN_455 = 5'h1d == fence_cnt ? d2_29 : _GEN_454; // @[DCache.scala 111:32 DCache.scala 111:32]
  wire  _GEN_456 = 5'h1e == fence_cnt ? d2_30 : _GEN_455; // @[DCache.scala 111:32 DCache.scala 111:32]
  wire  _GEN_457 = 5'h1f == fence_cnt ? d2_31 : _GEN_456; // @[DCache.scala 111:32 DCache.scala 111:32]
  wire [2:0] _GEN_458 = ~_GEN_457 | _GEN_457 & io_axi_wdone ? 3'h6 : state; // @[DCache.scala 111:91 DCache.scala 111:98 DCache.scala 69:24]
  wire  _T_17 = 3'h6 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_459 = _T_11 ? 3'h0 : 3'h5; // @[DCache.scala 114:54 DCache.scala 114:61 DCache.scala 115:31]
  wire [2:0] _GEN_460 = _T_17 ? _GEN_459 : state; // @[Conditional.scala 39:67 DCache.scala 69:24]
  wire [2:0] _GEN_461 = _T_12 ? _GEN_458 : _GEN_460; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_462 = _T_10 ? _GEN_425 : _GEN_461; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_463 = _T_5 ? _GEN_424 : _GEN_462; // @[Conditional.scala 39:67]
  wire  update = state == 3'h2 & io_axi_rvalid; // @[DCache.scala 121:39]
  wire  way1write = hit1 & op; // @[DCache.scala 122:26]
  wire  way2write = hit2 & op; // @[DCache.scala 123:26]
  wire  _T_19 = state == 3'h4; // @[DCache.scala 126:16]
  wire  _T_20 = update & updateway1; // @[DCache.scala 127:22]
  wire  _GEN_1182 = 5'h0 == index_addr; // @[DCache.scala 128:41 DCache.scala 128:41 DCache.scala 53:26]
  wire  _GEN_1183 = 5'h1 == index_addr; // @[DCache.scala 128:41 DCache.scala 128:41 DCache.scala 53:26]
  wire  _GEN_1184 = 5'h2 == index_addr; // @[DCache.scala 128:41 DCache.scala 128:41 DCache.scala 53:26]
  wire  _GEN_1185 = 5'h3 == index_addr; // @[DCache.scala 128:41 DCache.scala 128:41 DCache.scala 53:26]
  wire  _GEN_1186 = 5'h4 == index_addr; // @[DCache.scala 128:41 DCache.scala 128:41 DCache.scala 53:26]
  wire  _GEN_1187 = 5'h5 == index_addr; // @[DCache.scala 128:41 DCache.scala 128:41 DCache.scala 53:26]
  wire  _GEN_1188 = 5'h6 == index_addr; // @[DCache.scala 128:41 DCache.scala 128:41 DCache.scala 53:26]
  wire  _GEN_1189 = 5'h7 == index_addr; // @[DCache.scala 128:41 DCache.scala 128:41 DCache.scala 53:26]
  wire  _GEN_1190 = 5'h8 == index_addr; // @[DCache.scala 128:41 DCache.scala 128:41 DCache.scala 53:26]
  wire  _GEN_1191 = 5'h9 == index_addr; // @[DCache.scala 128:41 DCache.scala 128:41 DCache.scala 53:26]
  wire  _GEN_1192 = 5'ha == index_addr; // @[DCache.scala 128:41 DCache.scala 128:41 DCache.scala 53:26]
  wire  _GEN_1193 = 5'hb == index_addr; // @[DCache.scala 128:41 DCache.scala 128:41 DCache.scala 53:26]
  wire  _GEN_1194 = 5'hc == index_addr; // @[DCache.scala 128:41 DCache.scala 128:41 DCache.scala 53:26]
  wire  _GEN_1195 = 5'hd == index_addr; // @[DCache.scala 128:41 DCache.scala 128:41 DCache.scala 53:26]
  wire  _GEN_1196 = 5'he == index_addr; // @[DCache.scala 128:41 DCache.scala 128:41 DCache.scala 53:26]
  wire  _GEN_1197 = 5'hf == index_addr; // @[DCache.scala 128:41 DCache.scala 128:41 DCache.scala 53:26]
  wire  _GEN_1198 = 5'h10 == index_addr; // @[DCache.scala 128:41 DCache.scala 128:41 DCache.scala 53:26]
  wire  _GEN_1199 = 5'h11 == index_addr; // @[DCache.scala 128:41 DCache.scala 128:41 DCache.scala 53:26]
  wire  _GEN_1200 = 5'h12 == index_addr; // @[DCache.scala 128:41 DCache.scala 128:41 DCache.scala 53:26]
  wire  _GEN_1201 = 5'h13 == index_addr; // @[DCache.scala 128:41 DCache.scala 128:41 DCache.scala 53:26]
  wire  _GEN_1202 = 5'h14 == index_addr; // @[DCache.scala 128:41 DCache.scala 128:41 DCache.scala 53:26]
  wire  _GEN_1203 = 5'h15 == index_addr; // @[DCache.scala 128:41 DCache.scala 128:41 DCache.scala 53:26]
  wire  _GEN_1204 = 5'h16 == index_addr; // @[DCache.scala 128:41 DCache.scala 128:41 DCache.scala 53:26]
  wire  _GEN_1205 = 5'h17 == index_addr; // @[DCache.scala 128:41 DCache.scala 128:41 DCache.scala 53:26]
  wire  _GEN_1206 = 5'h18 == index_addr; // @[DCache.scala 128:41 DCache.scala 128:41 DCache.scala 53:26]
  wire  _GEN_1207 = 5'h19 == index_addr; // @[DCache.scala 128:41 DCache.scala 128:41 DCache.scala 53:26]
  wire  _GEN_1208 = 5'h1a == index_addr; // @[DCache.scala 128:41 DCache.scala 128:41 DCache.scala 53:26]
  wire  _GEN_1209 = 5'h1b == index_addr; // @[DCache.scala 128:41 DCache.scala 128:41 DCache.scala 53:26]
  wire  _GEN_1210 = 5'h1c == index_addr; // @[DCache.scala 128:41 DCache.scala 128:41 DCache.scala 53:26]
  wire  _GEN_1211 = 5'h1d == index_addr; // @[DCache.scala 128:41 DCache.scala 128:41 DCache.scala 53:26]
  wire  _GEN_1212 = 5'h1e == index_addr; // @[DCache.scala 128:41 DCache.scala 128:41 DCache.scala 53:26]
  wire  _GEN_1213 = 5'h1f == index_addr; // @[DCache.scala 128:41 DCache.scala 128:41 DCache.scala 53:26]
  wire  _T_21 = state == 3'h6; // @[DCache.scala 130:16]
  wire  _T_22 = update & updateway2; // @[DCache.scala 131:22]
  wire [7:0] mask64_hi_hi_hi_lo = wm[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] mask64_hi_hi_lo = wm[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] mask64_hi_lo_hi = wm[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] mask64_hi_lo_lo = wm[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] mask64_lo_hi_hi = wm[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] mask64_lo_hi_lo = wm[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] mask64_lo_lo_hi = wm[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] mask64_lo_lo_lo = wm[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [511:0] mask64 = {448'h0,mask64_hi_hi_hi_lo,mask64_hi_hi_lo,mask64_hi_lo_hi,mask64_hi_lo_lo,mask64_lo_hi_hi,
    mask64_lo_hi_lo,mask64_lo_lo_hi,mask64_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [8:0] _blockmask_T_1 = {offset_addr[5:3], 6'h0}; // @[DCache.scala 137:52]
  wire [1022:0] _GEN_1246 = {{511'd0}, mask64}; // @[DCache.scala 137:29]
  wire [1022:0] _blockmask_T_2 = _GEN_1246 << _blockmask_T_1; // @[DCache.scala 137:29]
  wire [511:0] blockmask = _blockmask_T_2[511:0]; // @[DCache.scala 137:58]
  wire [574:0] _GEN_1247 = {{511'd0}, wdata}; // @[DCache.scala 138:29]
  wire [574:0] _blockwdata_T_2 = _GEN_1247 << _blockmask_T_1; // @[DCache.scala 138:29]
  wire [511:0] blockwdata = _blockwdata_T_2[511:0]; // @[DCache.scala 138:58]
  wire [511:0] _block1_after_write_T = ~blockmask; // @[DCache.scala 139:53]
  wire [511:0] _block1_after_write_T_1 = _GEN_163 & _block1_after_write_T; // @[DCache.scala 139:50]
  wire [511:0] _block1_after_write_T_2 = blockmask & blockwdata; // @[DCache.scala 139:79]
  wire [511:0] block1_after_write = _block1_after_write_T_1 | _block1_after_write_T_2; // @[DCache.scala 139:66]
  wire [511:0] _block2_after_write_T_1 = _GEN_195 & _block1_after_write_T; // @[DCache.scala 140:50]
  wire [511:0] block2_after_write = _block2_after_write_T_1 | _block1_after_write_T_2; // @[DCache.scala 140:66]
  wire  _T_23 = state == 3'h3; // @[DCache.scala 157:16]
  wire [52:0] _GEN_1044 = 5'h1 == fence_cnt ? tag1_1 : tag1_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1045 = 5'h2 == fence_cnt ? tag1_2 : _GEN_1044; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1046 = 5'h3 == fence_cnt ? tag1_3 : _GEN_1045; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1047 = 5'h4 == fence_cnt ? tag1_4 : _GEN_1046; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1048 = 5'h5 == fence_cnt ? tag1_5 : _GEN_1047; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1049 = 5'h6 == fence_cnt ? tag1_6 : _GEN_1048; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1050 = 5'h7 == fence_cnt ? tag1_7 : _GEN_1049; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1051 = 5'h8 == fence_cnt ? tag1_8 : _GEN_1050; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1052 = 5'h9 == fence_cnt ? tag1_9 : _GEN_1051; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1053 = 5'ha == fence_cnt ? tag1_10 : _GEN_1052; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1054 = 5'hb == fence_cnt ? tag1_11 : _GEN_1053; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1055 = 5'hc == fence_cnt ? tag1_12 : _GEN_1054; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1056 = 5'hd == fence_cnt ? tag1_13 : _GEN_1055; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1057 = 5'he == fence_cnt ? tag1_14 : _GEN_1056; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1058 = 5'hf == fence_cnt ? tag1_15 : _GEN_1057; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1059 = 5'h10 == fence_cnt ? tag1_16 : _GEN_1058; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1060 = 5'h11 == fence_cnt ? tag1_17 : _GEN_1059; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1061 = 5'h12 == fence_cnt ? tag1_18 : _GEN_1060; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1062 = 5'h13 == fence_cnt ? tag1_19 : _GEN_1061; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1063 = 5'h14 == fence_cnt ? tag1_20 : _GEN_1062; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1064 = 5'h15 == fence_cnt ? tag1_21 : _GEN_1063; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1065 = 5'h16 == fence_cnt ? tag1_22 : _GEN_1064; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1066 = 5'h17 == fence_cnt ? tag1_23 : _GEN_1065; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1067 = 5'h18 == fence_cnt ? tag1_24 : _GEN_1066; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1068 = 5'h19 == fence_cnt ? tag1_25 : _GEN_1067; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1069 = 5'h1a == fence_cnt ? tag1_26 : _GEN_1068; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1070 = 5'h1b == fence_cnt ? tag1_27 : _GEN_1069; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1071 = 5'h1c == fence_cnt ? tag1_28 : _GEN_1070; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1072 = 5'h1d == fence_cnt ? tag1_29 : _GEN_1071; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1073 = 5'h1e == fence_cnt ? tag1_30 : _GEN_1072; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1074 = 5'h1f == fence_cnt ? tag1_31 : _GEN_1073; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [63:0] _io_axi_waddr_T = {_GEN_1074,fence_cnt,6'h0}; // @[Cat.scala 30:58]
  wire [511:0] _GEN_1076 = 5'h1 == fence_cnt ? block1_1 : block1_0; // @[DCache.scala 160:25 DCache.scala 160:25]
  wire [511:0] _GEN_1077 = 5'h2 == fence_cnt ? block1_2 : _GEN_1076; // @[DCache.scala 160:25 DCache.scala 160:25]
  wire [511:0] _GEN_1078 = 5'h3 == fence_cnt ? block1_3 : _GEN_1077; // @[DCache.scala 160:25 DCache.scala 160:25]
  wire [511:0] _GEN_1079 = 5'h4 == fence_cnt ? block1_4 : _GEN_1078; // @[DCache.scala 160:25 DCache.scala 160:25]
  wire [511:0] _GEN_1080 = 5'h5 == fence_cnt ? block1_5 : _GEN_1079; // @[DCache.scala 160:25 DCache.scala 160:25]
  wire [511:0] _GEN_1081 = 5'h6 == fence_cnt ? block1_6 : _GEN_1080; // @[DCache.scala 160:25 DCache.scala 160:25]
  wire [511:0] _GEN_1082 = 5'h7 == fence_cnt ? block1_7 : _GEN_1081; // @[DCache.scala 160:25 DCache.scala 160:25]
  wire [511:0] _GEN_1083 = 5'h8 == fence_cnt ? block1_8 : _GEN_1082; // @[DCache.scala 160:25 DCache.scala 160:25]
  wire [511:0] _GEN_1084 = 5'h9 == fence_cnt ? block1_9 : _GEN_1083; // @[DCache.scala 160:25 DCache.scala 160:25]
  wire [511:0] _GEN_1085 = 5'ha == fence_cnt ? block1_10 : _GEN_1084; // @[DCache.scala 160:25 DCache.scala 160:25]
  wire [511:0] _GEN_1086 = 5'hb == fence_cnt ? block1_11 : _GEN_1085; // @[DCache.scala 160:25 DCache.scala 160:25]
  wire [511:0] _GEN_1087 = 5'hc == fence_cnt ? block1_12 : _GEN_1086; // @[DCache.scala 160:25 DCache.scala 160:25]
  wire [511:0] _GEN_1088 = 5'hd == fence_cnt ? block1_13 : _GEN_1087; // @[DCache.scala 160:25 DCache.scala 160:25]
  wire [511:0] _GEN_1089 = 5'he == fence_cnt ? block1_14 : _GEN_1088; // @[DCache.scala 160:25 DCache.scala 160:25]
  wire [511:0] _GEN_1090 = 5'hf == fence_cnt ? block1_15 : _GEN_1089; // @[DCache.scala 160:25 DCache.scala 160:25]
  wire [511:0] _GEN_1091 = 5'h10 == fence_cnt ? block1_16 : _GEN_1090; // @[DCache.scala 160:25 DCache.scala 160:25]
  wire [511:0] _GEN_1092 = 5'h11 == fence_cnt ? block1_17 : _GEN_1091; // @[DCache.scala 160:25 DCache.scala 160:25]
  wire [511:0] _GEN_1093 = 5'h12 == fence_cnt ? block1_18 : _GEN_1092; // @[DCache.scala 160:25 DCache.scala 160:25]
  wire [511:0] _GEN_1094 = 5'h13 == fence_cnt ? block1_19 : _GEN_1093; // @[DCache.scala 160:25 DCache.scala 160:25]
  wire [511:0] _GEN_1095 = 5'h14 == fence_cnt ? block1_20 : _GEN_1094; // @[DCache.scala 160:25 DCache.scala 160:25]
  wire [511:0] _GEN_1096 = 5'h15 == fence_cnt ? block1_21 : _GEN_1095; // @[DCache.scala 160:25 DCache.scala 160:25]
  wire [511:0] _GEN_1097 = 5'h16 == fence_cnt ? block1_22 : _GEN_1096; // @[DCache.scala 160:25 DCache.scala 160:25]
  wire [511:0] _GEN_1098 = 5'h17 == fence_cnt ? block1_23 : _GEN_1097; // @[DCache.scala 160:25 DCache.scala 160:25]
  wire [511:0] _GEN_1099 = 5'h18 == fence_cnt ? block1_24 : _GEN_1098; // @[DCache.scala 160:25 DCache.scala 160:25]
  wire [511:0] _GEN_1100 = 5'h19 == fence_cnt ? block1_25 : _GEN_1099; // @[DCache.scala 160:25 DCache.scala 160:25]
  wire [511:0] _GEN_1101 = 5'h1a == fence_cnt ? block1_26 : _GEN_1100; // @[DCache.scala 160:25 DCache.scala 160:25]
  wire [511:0] _GEN_1102 = 5'h1b == fence_cnt ? block1_27 : _GEN_1101; // @[DCache.scala 160:25 DCache.scala 160:25]
  wire [511:0] _GEN_1103 = 5'h1c == fence_cnt ? block1_28 : _GEN_1102; // @[DCache.scala 160:25 DCache.scala 160:25]
  wire [511:0] _GEN_1104 = 5'h1d == fence_cnt ? block1_29 : _GEN_1103; // @[DCache.scala 160:25 DCache.scala 160:25]
  wire [511:0] _GEN_1105 = 5'h1e == fence_cnt ? block1_30 : _GEN_1104; // @[DCache.scala 160:25 DCache.scala 160:25]
  wire [511:0] _GEN_1106 = 5'h1f == fence_cnt ? block1_31 : _GEN_1105; // @[DCache.scala 160:25 DCache.scala 160:25]
  wire  _T_25 = state == 3'h5; // @[DCache.scala 162:21]
  wire [52:0] _GEN_1108 = 5'h1 == fence_cnt ? tag2_1 : tag2_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1109 = 5'h2 == fence_cnt ? tag2_2 : _GEN_1108; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1110 = 5'h3 == fence_cnt ? tag2_3 : _GEN_1109; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1111 = 5'h4 == fence_cnt ? tag2_4 : _GEN_1110; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1112 = 5'h5 == fence_cnt ? tag2_5 : _GEN_1111; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1113 = 5'h6 == fence_cnt ? tag2_6 : _GEN_1112; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1114 = 5'h7 == fence_cnt ? tag2_7 : _GEN_1113; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1115 = 5'h8 == fence_cnt ? tag2_8 : _GEN_1114; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1116 = 5'h9 == fence_cnt ? tag2_9 : _GEN_1115; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1117 = 5'ha == fence_cnt ? tag2_10 : _GEN_1116; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1118 = 5'hb == fence_cnt ? tag2_11 : _GEN_1117; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1119 = 5'hc == fence_cnt ? tag2_12 : _GEN_1118; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1120 = 5'hd == fence_cnt ? tag2_13 : _GEN_1119; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1121 = 5'he == fence_cnt ? tag2_14 : _GEN_1120; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1122 = 5'hf == fence_cnt ? tag2_15 : _GEN_1121; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1123 = 5'h10 == fence_cnt ? tag2_16 : _GEN_1122; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1124 = 5'h11 == fence_cnt ? tag2_17 : _GEN_1123; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1125 = 5'h12 == fence_cnt ? tag2_18 : _GEN_1124; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1126 = 5'h13 == fence_cnt ? tag2_19 : _GEN_1125; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1127 = 5'h14 == fence_cnt ? tag2_20 : _GEN_1126; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1128 = 5'h15 == fence_cnt ? tag2_21 : _GEN_1127; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1129 = 5'h16 == fence_cnt ? tag2_22 : _GEN_1128; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1130 = 5'h17 == fence_cnt ? tag2_23 : _GEN_1129; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1131 = 5'h18 == fence_cnt ? tag2_24 : _GEN_1130; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1132 = 5'h19 == fence_cnt ? tag2_25 : _GEN_1131; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1133 = 5'h1a == fence_cnt ? tag2_26 : _GEN_1132; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1134 = 5'h1b == fence_cnt ? tag2_27 : _GEN_1133; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1135 = 5'h1c == fence_cnt ? tag2_28 : _GEN_1134; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1136 = 5'h1d == fence_cnt ? tag2_29 : _GEN_1135; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1137 = 5'h1e == fence_cnt ? tag2_30 : _GEN_1136; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [52:0] _GEN_1138 = 5'h1f == fence_cnt ? tag2_31 : _GEN_1137; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [63:0] _io_axi_waddr_T_1 = {_GEN_1138,fence_cnt,6'h0}; // @[Cat.scala 30:58]
  wire [511:0] _GEN_1140 = 5'h1 == fence_cnt ? block2_1 : block2_0; // @[DCache.scala 165:25 DCache.scala 165:25]
  wire [511:0] _GEN_1141 = 5'h2 == fence_cnt ? block2_2 : _GEN_1140; // @[DCache.scala 165:25 DCache.scala 165:25]
  wire [511:0] _GEN_1142 = 5'h3 == fence_cnt ? block2_3 : _GEN_1141; // @[DCache.scala 165:25 DCache.scala 165:25]
  wire [511:0] _GEN_1143 = 5'h4 == fence_cnt ? block2_4 : _GEN_1142; // @[DCache.scala 165:25 DCache.scala 165:25]
  wire [511:0] _GEN_1144 = 5'h5 == fence_cnt ? block2_5 : _GEN_1143; // @[DCache.scala 165:25 DCache.scala 165:25]
  wire [511:0] _GEN_1145 = 5'h6 == fence_cnt ? block2_6 : _GEN_1144; // @[DCache.scala 165:25 DCache.scala 165:25]
  wire [511:0] _GEN_1146 = 5'h7 == fence_cnt ? block2_7 : _GEN_1145; // @[DCache.scala 165:25 DCache.scala 165:25]
  wire [511:0] _GEN_1147 = 5'h8 == fence_cnt ? block2_8 : _GEN_1146; // @[DCache.scala 165:25 DCache.scala 165:25]
  wire [511:0] _GEN_1148 = 5'h9 == fence_cnt ? block2_9 : _GEN_1147; // @[DCache.scala 165:25 DCache.scala 165:25]
  wire [511:0] _GEN_1149 = 5'ha == fence_cnt ? block2_10 : _GEN_1148; // @[DCache.scala 165:25 DCache.scala 165:25]
  wire [511:0] _GEN_1150 = 5'hb == fence_cnt ? block2_11 : _GEN_1149; // @[DCache.scala 165:25 DCache.scala 165:25]
  wire [511:0] _GEN_1151 = 5'hc == fence_cnt ? block2_12 : _GEN_1150; // @[DCache.scala 165:25 DCache.scala 165:25]
  wire [511:0] _GEN_1152 = 5'hd == fence_cnt ? block2_13 : _GEN_1151; // @[DCache.scala 165:25 DCache.scala 165:25]
  wire [511:0] _GEN_1153 = 5'he == fence_cnt ? block2_14 : _GEN_1152; // @[DCache.scala 165:25 DCache.scala 165:25]
  wire [511:0] _GEN_1154 = 5'hf == fence_cnt ? block2_15 : _GEN_1153; // @[DCache.scala 165:25 DCache.scala 165:25]
  wire [511:0] _GEN_1155 = 5'h10 == fence_cnt ? block2_16 : _GEN_1154; // @[DCache.scala 165:25 DCache.scala 165:25]
  wire [511:0] _GEN_1156 = 5'h11 == fence_cnt ? block2_17 : _GEN_1155; // @[DCache.scala 165:25 DCache.scala 165:25]
  wire [511:0] _GEN_1157 = 5'h12 == fence_cnt ? block2_18 : _GEN_1156; // @[DCache.scala 165:25 DCache.scala 165:25]
  wire [511:0] _GEN_1158 = 5'h13 == fence_cnt ? block2_19 : _GEN_1157; // @[DCache.scala 165:25 DCache.scala 165:25]
  wire [511:0] _GEN_1159 = 5'h14 == fence_cnt ? block2_20 : _GEN_1158; // @[DCache.scala 165:25 DCache.scala 165:25]
  wire [511:0] _GEN_1160 = 5'h15 == fence_cnt ? block2_21 : _GEN_1159; // @[DCache.scala 165:25 DCache.scala 165:25]
  wire [511:0] _GEN_1161 = 5'h16 == fence_cnt ? block2_22 : _GEN_1160; // @[DCache.scala 165:25 DCache.scala 165:25]
  wire [511:0] _GEN_1162 = 5'h17 == fence_cnt ? block2_23 : _GEN_1161; // @[DCache.scala 165:25 DCache.scala 165:25]
  wire [511:0] _GEN_1163 = 5'h18 == fence_cnt ? block2_24 : _GEN_1162; // @[DCache.scala 165:25 DCache.scala 165:25]
  wire [511:0] _GEN_1164 = 5'h19 == fence_cnt ? block2_25 : _GEN_1163; // @[DCache.scala 165:25 DCache.scala 165:25]
  wire [511:0] _GEN_1165 = 5'h1a == fence_cnt ? block2_26 : _GEN_1164; // @[DCache.scala 165:25 DCache.scala 165:25]
  wire [511:0] _GEN_1166 = 5'h1b == fence_cnt ? block2_27 : _GEN_1165; // @[DCache.scala 165:25 DCache.scala 165:25]
  wire [511:0] _GEN_1167 = 5'h1c == fence_cnt ? block2_28 : _GEN_1166; // @[DCache.scala 165:25 DCache.scala 165:25]
  wire [511:0] _GEN_1168 = 5'h1d == fence_cnt ? block2_29 : _GEN_1167; // @[DCache.scala 165:25 DCache.scala 165:25]
  wire [511:0] _GEN_1169 = 5'h1e == fence_cnt ? block2_30 : _GEN_1168; // @[DCache.scala 165:25 DCache.scala 165:25]
  wire [511:0] _GEN_1170 = 5'h1f == fence_cnt ? block2_31 : _GEN_1169; // @[DCache.scala 165:25 DCache.scala 165:25]
  wire [52:0] io_axi_waddr_hi_hi = updateway1 ? _GEN_35 : _GEN_99; // @[DCache.scala 169:35]
  wire [63:0] _io_axi_waddr_T_2 = {io_axi_waddr_hi_hi,index_addr,6'h0}; // @[Cat.scala 30:58]
  wire [511:0] _io_axi_wdata_T = updateway1 ? _GEN_163 : _GEN_195; // @[DCache.scala 170:31]
  wire  _GEN_1171 = state == 3'h1 & state == 3'h1; // @[DCache.scala 167:36 DCache.scala 168:25 DCache.scala 173:25]
  wire [63:0] _GEN_1172 = state == 3'h1 ? _io_axi_waddr_T_2 : 64'h0; // @[DCache.scala 167:36 DCache.scala 169:25 DCache.scala 174:25]
  wire [511:0] _GEN_1173 = state == 3'h1 ? _io_axi_wdata_T : 512'h0; // @[DCache.scala 167:36 DCache.scala 170:25 DCache.scala 175:25]
  wire  _GEN_1174 = state == 3'h5 & _GEN_457 | _GEN_1171; // @[DCache.scala 162:55 DCache.scala 163:25]
  wire [63:0] _GEN_1175 = state == 3'h5 & _GEN_457 ? _io_axi_waddr_T_1 : _GEN_1172; // @[DCache.scala 162:55 DCache.scala 164:25]
  wire [511:0] _GEN_1176 = state == 3'h5 & _GEN_457 ? _GEN_1170 : _GEN_1173; // @[DCache.scala 162:55 DCache.scala 165:25]
  wire [4:0] _lo_T_1 = fence_cnt + 5'h1; // @[DCache.scala 180:87]
  assign io_dmem_ok = (hit | not_en_yet) & state == 3'h0; // @[DCache.scala 78:44]
  assign io_dmem_rdata = hit2 ? rdata2 : _rdata_T; // @[DCache.scala 72:26]
  assign io_axi_req = state == 3'h2; // @[DCache.scala 151:30]
  assign io_axi_raddr = addr & 64'hffffffffffffffc0; // @[DCache.scala 152:29]
  assign io_axi_weq = state == 3'h3 & _GEN_423 | _GEN_1174; // @[DCache.scala 157:50 DCache.scala 158:25]
  assign io_axi_waddr = state == 3'h3 & _GEN_423 ? _io_axi_waddr_T : _GEN_1175; // @[DCache.scala 157:50 DCache.scala 159:25]
  assign io_axi_wdata = state == 3'h3 & _GEN_423 ? _GEN_1106 : _GEN_1176; // @[DCache.scala 157:50 DCache.scala 160:25]
  assign io_fence_done = _T_21 & _T_11; // @[DCache.scala 185:47]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 27:20]
      op <= 1'h0; // @[Reg.scala 27:20]
    end else if (_op_T) begin // @[Reg.scala 28:19]
      op <= io_dmem_op; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      addr <= 64'h0; // @[Reg.scala 27:20]
    end else if (_op_T) begin // @[Reg.scala 28:19]
      addr <= _addr_T; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      wdata <= 64'h0; // @[Reg.scala 27:20]
    end else if (_op_T) begin // @[Reg.scala 28:19]
      wdata <= io_dmem_wdata; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      wm <= 8'h0; // @[Reg.scala 27:20]
    end else if (_op_T) begin // @[Reg.scala 28:19]
      wm <= io_dmem_wmask; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[DCache.scala 52:26]
      v1_0 <= 1'h0; // @[DCache.scala 52:26]
    end else if (5'h0 == index_addr) begin // @[DCache.scala 145:26]
      v1_0 <= _T_20 | _GEN_67; // @[DCache.scala 145:26]
    end
    if (reset) begin // @[DCache.scala 52:26]
      v1_1 <= 1'h0; // @[DCache.scala 52:26]
    end else if (5'h1 == index_addr) begin // @[DCache.scala 145:26]
      v1_1 <= _T_20 | _GEN_67; // @[DCache.scala 145:26]
    end
    if (reset) begin // @[DCache.scala 52:26]
      v1_2 <= 1'h0; // @[DCache.scala 52:26]
    end else if (5'h2 == index_addr) begin // @[DCache.scala 145:26]
      v1_2 <= _T_20 | _GEN_67; // @[DCache.scala 145:26]
    end
    if (reset) begin // @[DCache.scala 52:26]
      v1_3 <= 1'h0; // @[DCache.scala 52:26]
    end else if (5'h3 == index_addr) begin // @[DCache.scala 145:26]
      v1_3 <= _T_20 | _GEN_67; // @[DCache.scala 145:26]
    end
    if (reset) begin // @[DCache.scala 52:26]
      v1_4 <= 1'h0; // @[DCache.scala 52:26]
    end else if (5'h4 == index_addr) begin // @[DCache.scala 145:26]
      v1_4 <= _T_20 | _GEN_67; // @[DCache.scala 145:26]
    end
    if (reset) begin // @[DCache.scala 52:26]
      v1_5 <= 1'h0; // @[DCache.scala 52:26]
    end else if (5'h5 == index_addr) begin // @[DCache.scala 145:26]
      v1_5 <= _T_20 | _GEN_67; // @[DCache.scala 145:26]
    end
    if (reset) begin // @[DCache.scala 52:26]
      v1_6 <= 1'h0; // @[DCache.scala 52:26]
    end else if (5'h6 == index_addr) begin // @[DCache.scala 145:26]
      v1_6 <= _T_20 | _GEN_67; // @[DCache.scala 145:26]
    end
    if (reset) begin // @[DCache.scala 52:26]
      v1_7 <= 1'h0; // @[DCache.scala 52:26]
    end else if (5'h7 == index_addr) begin // @[DCache.scala 145:26]
      v1_7 <= _T_20 | _GEN_67; // @[DCache.scala 145:26]
    end
    if (reset) begin // @[DCache.scala 52:26]
      v1_8 <= 1'h0; // @[DCache.scala 52:26]
    end else if (5'h8 == index_addr) begin // @[DCache.scala 145:26]
      v1_8 <= _T_20 | _GEN_67; // @[DCache.scala 145:26]
    end
    if (reset) begin // @[DCache.scala 52:26]
      v1_9 <= 1'h0; // @[DCache.scala 52:26]
    end else if (5'h9 == index_addr) begin // @[DCache.scala 145:26]
      v1_9 <= _T_20 | _GEN_67; // @[DCache.scala 145:26]
    end
    if (reset) begin // @[DCache.scala 52:26]
      v1_10 <= 1'h0; // @[DCache.scala 52:26]
    end else if (5'ha == index_addr) begin // @[DCache.scala 145:26]
      v1_10 <= _T_20 | _GEN_67; // @[DCache.scala 145:26]
    end
    if (reset) begin // @[DCache.scala 52:26]
      v1_11 <= 1'h0; // @[DCache.scala 52:26]
    end else if (5'hb == index_addr) begin // @[DCache.scala 145:26]
      v1_11 <= _T_20 | _GEN_67; // @[DCache.scala 145:26]
    end
    if (reset) begin // @[DCache.scala 52:26]
      v1_12 <= 1'h0; // @[DCache.scala 52:26]
    end else if (5'hc == index_addr) begin // @[DCache.scala 145:26]
      v1_12 <= _T_20 | _GEN_67; // @[DCache.scala 145:26]
    end
    if (reset) begin // @[DCache.scala 52:26]
      v1_13 <= 1'h0; // @[DCache.scala 52:26]
    end else if (5'hd == index_addr) begin // @[DCache.scala 145:26]
      v1_13 <= _T_20 | _GEN_67; // @[DCache.scala 145:26]
    end
    if (reset) begin // @[DCache.scala 52:26]
      v1_14 <= 1'h0; // @[DCache.scala 52:26]
    end else if (5'he == index_addr) begin // @[DCache.scala 145:26]
      v1_14 <= _T_20 | _GEN_67; // @[DCache.scala 145:26]
    end
    if (reset) begin // @[DCache.scala 52:26]
      v1_15 <= 1'h0; // @[DCache.scala 52:26]
    end else if (5'hf == index_addr) begin // @[DCache.scala 145:26]
      v1_15 <= _T_20 | _GEN_67; // @[DCache.scala 145:26]
    end
    if (reset) begin // @[DCache.scala 52:26]
      v1_16 <= 1'h0; // @[DCache.scala 52:26]
    end else if (5'h10 == index_addr) begin // @[DCache.scala 145:26]
      v1_16 <= _T_20 | _GEN_67; // @[DCache.scala 145:26]
    end
    if (reset) begin // @[DCache.scala 52:26]
      v1_17 <= 1'h0; // @[DCache.scala 52:26]
    end else if (5'h11 == index_addr) begin // @[DCache.scala 145:26]
      v1_17 <= _T_20 | _GEN_67; // @[DCache.scala 145:26]
    end
    if (reset) begin // @[DCache.scala 52:26]
      v1_18 <= 1'h0; // @[DCache.scala 52:26]
    end else if (5'h12 == index_addr) begin // @[DCache.scala 145:26]
      v1_18 <= _T_20 | _GEN_67; // @[DCache.scala 145:26]
    end
    if (reset) begin // @[DCache.scala 52:26]
      v1_19 <= 1'h0; // @[DCache.scala 52:26]
    end else if (5'h13 == index_addr) begin // @[DCache.scala 145:26]
      v1_19 <= _T_20 | _GEN_67; // @[DCache.scala 145:26]
    end
    if (reset) begin // @[DCache.scala 52:26]
      v1_20 <= 1'h0; // @[DCache.scala 52:26]
    end else if (5'h14 == index_addr) begin // @[DCache.scala 145:26]
      v1_20 <= _T_20 | _GEN_67; // @[DCache.scala 145:26]
    end
    if (reset) begin // @[DCache.scala 52:26]
      v1_21 <= 1'h0; // @[DCache.scala 52:26]
    end else if (5'h15 == index_addr) begin // @[DCache.scala 145:26]
      v1_21 <= _T_20 | _GEN_67; // @[DCache.scala 145:26]
    end
    if (reset) begin // @[DCache.scala 52:26]
      v1_22 <= 1'h0; // @[DCache.scala 52:26]
    end else if (5'h16 == index_addr) begin // @[DCache.scala 145:26]
      v1_22 <= _T_20 | _GEN_67; // @[DCache.scala 145:26]
    end
    if (reset) begin // @[DCache.scala 52:26]
      v1_23 <= 1'h0; // @[DCache.scala 52:26]
    end else if (5'h17 == index_addr) begin // @[DCache.scala 145:26]
      v1_23 <= _T_20 | _GEN_67; // @[DCache.scala 145:26]
    end
    if (reset) begin // @[DCache.scala 52:26]
      v1_24 <= 1'h0; // @[DCache.scala 52:26]
    end else if (5'h18 == index_addr) begin // @[DCache.scala 145:26]
      v1_24 <= _T_20 | _GEN_67; // @[DCache.scala 145:26]
    end
    if (reset) begin // @[DCache.scala 52:26]
      v1_25 <= 1'h0; // @[DCache.scala 52:26]
    end else if (5'h19 == index_addr) begin // @[DCache.scala 145:26]
      v1_25 <= _T_20 | _GEN_67; // @[DCache.scala 145:26]
    end
    if (reset) begin // @[DCache.scala 52:26]
      v1_26 <= 1'h0; // @[DCache.scala 52:26]
    end else if (5'h1a == index_addr) begin // @[DCache.scala 145:26]
      v1_26 <= _T_20 | _GEN_67; // @[DCache.scala 145:26]
    end
    if (reset) begin // @[DCache.scala 52:26]
      v1_27 <= 1'h0; // @[DCache.scala 52:26]
    end else if (5'h1b == index_addr) begin // @[DCache.scala 145:26]
      v1_27 <= _T_20 | _GEN_67; // @[DCache.scala 145:26]
    end
    if (reset) begin // @[DCache.scala 52:26]
      v1_28 <= 1'h0; // @[DCache.scala 52:26]
    end else if (5'h1c == index_addr) begin // @[DCache.scala 145:26]
      v1_28 <= _T_20 | _GEN_67; // @[DCache.scala 145:26]
    end
    if (reset) begin // @[DCache.scala 52:26]
      v1_29 <= 1'h0; // @[DCache.scala 52:26]
    end else if (5'h1d == index_addr) begin // @[DCache.scala 145:26]
      v1_29 <= _T_20 | _GEN_67; // @[DCache.scala 145:26]
    end
    if (reset) begin // @[DCache.scala 52:26]
      v1_30 <= 1'h0; // @[DCache.scala 52:26]
    end else if (5'h1e == index_addr) begin // @[DCache.scala 145:26]
      v1_30 <= _T_20 | _GEN_67; // @[DCache.scala 145:26]
    end
    if (reset) begin // @[DCache.scala 52:26]
      v1_31 <= 1'h0; // @[DCache.scala 52:26]
    end else if (5'h1f == index_addr) begin // @[DCache.scala 145:26]
      v1_31 <= _T_20 | _GEN_67; // @[DCache.scala 145:26]
    end
    if (reset) begin // @[DCache.scala 53:26]
      d1_0 <= 1'h0; // @[DCache.scala 53:26]
    end else if (state == 3'h4) begin // @[DCache.scala 126:35]
      if (5'h0 == fence_cnt) begin // @[DCache.scala 126:50]
        d1_0 <= 1'h0; // @[DCache.scala 126:50]
      end
    end else if (update & updateway1) begin // @[DCache.scala 127:36]
      if (5'h0 == index_addr) begin // @[DCache.scala 127:52]
        d1_0 <= 1'h0; // @[DCache.scala 127:52]
      end
    end else if (way1write) begin // @[DCache.scala 128:25]
      d1_0 <= 5'h0 == index_addr | d1_0;
    end
    if (reset) begin // @[DCache.scala 53:26]
      d1_1 <= 1'h0; // @[DCache.scala 53:26]
    end else if (state == 3'h4) begin // @[DCache.scala 126:35]
      if (5'h1 == fence_cnt) begin // @[DCache.scala 126:50]
        d1_1 <= 1'h0; // @[DCache.scala 126:50]
      end
    end else if (update & updateway1) begin // @[DCache.scala 127:36]
      if (5'h1 == index_addr) begin // @[DCache.scala 127:52]
        d1_1 <= 1'h0; // @[DCache.scala 127:52]
      end
    end else if (way1write) begin // @[DCache.scala 128:25]
      d1_1 <= 5'h1 == index_addr | d1_1;
    end
    if (reset) begin // @[DCache.scala 53:26]
      d1_2 <= 1'h0; // @[DCache.scala 53:26]
    end else if (state == 3'h4) begin // @[DCache.scala 126:35]
      if (5'h2 == fence_cnt) begin // @[DCache.scala 126:50]
        d1_2 <= 1'h0; // @[DCache.scala 126:50]
      end
    end else if (update & updateway1) begin // @[DCache.scala 127:36]
      if (5'h2 == index_addr) begin // @[DCache.scala 127:52]
        d1_2 <= 1'h0; // @[DCache.scala 127:52]
      end
    end else if (way1write) begin // @[DCache.scala 128:25]
      d1_2 <= 5'h2 == index_addr | d1_2;
    end
    if (reset) begin // @[DCache.scala 53:26]
      d1_3 <= 1'h0; // @[DCache.scala 53:26]
    end else if (state == 3'h4) begin // @[DCache.scala 126:35]
      if (5'h3 == fence_cnt) begin // @[DCache.scala 126:50]
        d1_3 <= 1'h0; // @[DCache.scala 126:50]
      end
    end else if (update & updateway1) begin // @[DCache.scala 127:36]
      if (5'h3 == index_addr) begin // @[DCache.scala 127:52]
        d1_3 <= 1'h0; // @[DCache.scala 127:52]
      end
    end else if (way1write) begin // @[DCache.scala 128:25]
      d1_3 <= 5'h3 == index_addr | d1_3;
    end
    if (reset) begin // @[DCache.scala 53:26]
      d1_4 <= 1'h0; // @[DCache.scala 53:26]
    end else if (state == 3'h4) begin // @[DCache.scala 126:35]
      if (5'h4 == fence_cnt) begin // @[DCache.scala 126:50]
        d1_4 <= 1'h0; // @[DCache.scala 126:50]
      end
    end else if (update & updateway1) begin // @[DCache.scala 127:36]
      if (5'h4 == index_addr) begin // @[DCache.scala 127:52]
        d1_4 <= 1'h0; // @[DCache.scala 127:52]
      end
    end else if (way1write) begin // @[DCache.scala 128:25]
      d1_4 <= 5'h4 == index_addr | d1_4;
    end
    if (reset) begin // @[DCache.scala 53:26]
      d1_5 <= 1'h0; // @[DCache.scala 53:26]
    end else if (state == 3'h4) begin // @[DCache.scala 126:35]
      if (5'h5 == fence_cnt) begin // @[DCache.scala 126:50]
        d1_5 <= 1'h0; // @[DCache.scala 126:50]
      end
    end else if (update & updateway1) begin // @[DCache.scala 127:36]
      if (5'h5 == index_addr) begin // @[DCache.scala 127:52]
        d1_5 <= 1'h0; // @[DCache.scala 127:52]
      end
    end else if (way1write) begin // @[DCache.scala 128:25]
      d1_5 <= 5'h5 == index_addr | d1_5;
    end
    if (reset) begin // @[DCache.scala 53:26]
      d1_6 <= 1'h0; // @[DCache.scala 53:26]
    end else if (state == 3'h4) begin // @[DCache.scala 126:35]
      if (5'h6 == fence_cnt) begin // @[DCache.scala 126:50]
        d1_6 <= 1'h0; // @[DCache.scala 126:50]
      end
    end else if (update & updateway1) begin // @[DCache.scala 127:36]
      if (5'h6 == index_addr) begin // @[DCache.scala 127:52]
        d1_6 <= 1'h0; // @[DCache.scala 127:52]
      end
    end else if (way1write) begin // @[DCache.scala 128:25]
      d1_6 <= 5'h6 == index_addr | d1_6;
    end
    if (reset) begin // @[DCache.scala 53:26]
      d1_7 <= 1'h0; // @[DCache.scala 53:26]
    end else if (state == 3'h4) begin // @[DCache.scala 126:35]
      if (5'h7 == fence_cnt) begin // @[DCache.scala 126:50]
        d1_7 <= 1'h0; // @[DCache.scala 126:50]
      end
    end else if (update & updateway1) begin // @[DCache.scala 127:36]
      if (5'h7 == index_addr) begin // @[DCache.scala 127:52]
        d1_7 <= 1'h0; // @[DCache.scala 127:52]
      end
    end else if (way1write) begin // @[DCache.scala 128:25]
      d1_7 <= 5'h7 == index_addr | d1_7;
    end
    if (reset) begin // @[DCache.scala 53:26]
      d1_8 <= 1'h0; // @[DCache.scala 53:26]
    end else if (state == 3'h4) begin // @[DCache.scala 126:35]
      if (5'h8 == fence_cnt) begin // @[DCache.scala 126:50]
        d1_8 <= 1'h0; // @[DCache.scala 126:50]
      end
    end else if (update & updateway1) begin // @[DCache.scala 127:36]
      if (5'h8 == index_addr) begin // @[DCache.scala 127:52]
        d1_8 <= 1'h0; // @[DCache.scala 127:52]
      end
    end else if (way1write) begin // @[DCache.scala 128:25]
      d1_8 <= 5'h8 == index_addr | d1_8;
    end
    if (reset) begin // @[DCache.scala 53:26]
      d1_9 <= 1'h0; // @[DCache.scala 53:26]
    end else if (state == 3'h4) begin // @[DCache.scala 126:35]
      if (5'h9 == fence_cnt) begin // @[DCache.scala 126:50]
        d1_9 <= 1'h0; // @[DCache.scala 126:50]
      end
    end else if (update & updateway1) begin // @[DCache.scala 127:36]
      if (5'h9 == index_addr) begin // @[DCache.scala 127:52]
        d1_9 <= 1'h0; // @[DCache.scala 127:52]
      end
    end else if (way1write) begin // @[DCache.scala 128:25]
      d1_9 <= 5'h9 == index_addr | d1_9;
    end
    if (reset) begin // @[DCache.scala 53:26]
      d1_10 <= 1'h0; // @[DCache.scala 53:26]
    end else if (state == 3'h4) begin // @[DCache.scala 126:35]
      if (5'ha == fence_cnt) begin // @[DCache.scala 126:50]
        d1_10 <= 1'h0; // @[DCache.scala 126:50]
      end
    end else if (update & updateway1) begin // @[DCache.scala 127:36]
      if (5'ha == index_addr) begin // @[DCache.scala 127:52]
        d1_10 <= 1'h0; // @[DCache.scala 127:52]
      end
    end else if (way1write) begin // @[DCache.scala 128:25]
      d1_10 <= 5'ha == index_addr | d1_10;
    end
    if (reset) begin // @[DCache.scala 53:26]
      d1_11 <= 1'h0; // @[DCache.scala 53:26]
    end else if (state == 3'h4) begin // @[DCache.scala 126:35]
      if (5'hb == fence_cnt) begin // @[DCache.scala 126:50]
        d1_11 <= 1'h0; // @[DCache.scala 126:50]
      end
    end else if (update & updateway1) begin // @[DCache.scala 127:36]
      if (5'hb == index_addr) begin // @[DCache.scala 127:52]
        d1_11 <= 1'h0; // @[DCache.scala 127:52]
      end
    end else if (way1write) begin // @[DCache.scala 128:25]
      d1_11 <= 5'hb == index_addr | d1_11;
    end
    if (reset) begin // @[DCache.scala 53:26]
      d1_12 <= 1'h0; // @[DCache.scala 53:26]
    end else if (state == 3'h4) begin // @[DCache.scala 126:35]
      if (5'hc == fence_cnt) begin // @[DCache.scala 126:50]
        d1_12 <= 1'h0; // @[DCache.scala 126:50]
      end
    end else if (update & updateway1) begin // @[DCache.scala 127:36]
      if (5'hc == index_addr) begin // @[DCache.scala 127:52]
        d1_12 <= 1'h0; // @[DCache.scala 127:52]
      end
    end else if (way1write) begin // @[DCache.scala 128:25]
      d1_12 <= 5'hc == index_addr | d1_12;
    end
    if (reset) begin // @[DCache.scala 53:26]
      d1_13 <= 1'h0; // @[DCache.scala 53:26]
    end else if (state == 3'h4) begin // @[DCache.scala 126:35]
      if (5'hd == fence_cnt) begin // @[DCache.scala 126:50]
        d1_13 <= 1'h0; // @[DCache.scala 126:50]
      end
    end else if (update & updateway1) begin // @[DCache.scala 127:36]
      if (5'hd == index_addr) begin // @[DCache.scala 127:52]
        d1_13 <= 1'h0; // @[DCache.scala 127:52]
      end
    end else if (way1write) begin // @[DCache.scala 128:25]
      d1_13 <= 5'hd == index_addr | d1_13;
    end
    if (reset) begin // @[DCache.scala 53:26]
      d1_14 <= 1'h0; // @[DCache.scala 53:26]
    end else if (state == 3'h4) begin // @[DCache.scala 126:35]
      if (5'he == fence_cnt) begin // @[DCache.scala 126:50]
        d1_14 <= 1'h0; // @[DCache.scala 126:50]
      end
    end else if (update & updateway1) begin // @[DCache.scala 127:36]
      if (5'he == index_addr) begin // @[DCache.scala 127:52]
        d1_14 <= 1'h0; // @[DCache.scala 127:52]
      end
    end else if (way1write) begin // @[DCache.scala 128:25]
      d1_14 <= 5'he == index_addr | d1_14;
    end
    if (reset) begin // @[DCache.scala 53:26]
      d1_15 <= 1'h0; // @[DCache.scala 53:26]
    end else if (state == 3'h4) begin // @[DCache.scala 126:35]
      if (5'hf == fence_cnt) begin // @[DCache.scala 126:50]
        d1_15 <= 1'h0; // @[DCache.scala 126:50]
      end
    end else if (update & updateway1) begin // @[DCache.scala 127:36]
      if (5'hf == index_addr) begin // @[DCache.scala 127:52]
        d1_15 <= 1'h0; // @[DCache.scala 127:52]
      end
    end else if (way1write) begin // @[DCache.scala 128:25]
      d1_15 <= 5'hf == index_addr | d1_15;
    end
    if (reset) begin // @[DCache.scala 53:26]
      d1_16 <= 1'h0; // @[DCache.scala 53:26]
    end else if (state == 3'h4) begin // @[DCache.scala 126:35]
      if (5'h10 == fence_cnt) begin // @[DCache.scala 126:50]
        d1_16 <= 1'h0; // @[DCache.scala 126:50]
      end
    end else if (update & updateway1) begin // @[DCache.scala 127:36]
      if (5'h10 == index_addr) begin // @[DCache.scala 127:52]
        d1_16 <= 1'h0; // @[DCache.scala 127:52]
      end
    end else if (way1write) begin // @[DCache.scala 128:25]
      d1_16 <= 5'h10 == index_addr | d1_16;
    end
    if (reset) begin // @[DCache.scala 53:26]
      d1_17 <= 1'h0; // @[DCache.scala 53:26]
    end else if (state == 3'h4) begin // @[DCache.scala 126:35]
      if (5'h11 == fence_cnt) begin // @[DCache.scala 126:50]
        d1_17 <= 1'h0; // @[DCache.scala 126:50]
      end
    end else if (update & updateway1) begin // @[DCache.scala 127:36]
      if (5'h11 == index_addr) begin // @[DCache.scala 127:52]
        d1_17 <= 1'h0; // @[DCache.scala 127:52]
      end
    end else if (way1write) begin // @[DCache.scala 128:25]
      d1_17 <= 5'h11 == index_addr | d1_17;
    end
    if (reset) begin // @[DCache.scala 53:26]
      d1_18 <= 1'h0; // @[DCache.scala 53:26]
    end else if (state == 3'h4) begin // @[DCache.scala 126:35]
      if (5'h12 == fence_cnt) begin // @[DCache.scala 126:50]
        d1_18 <= 1'h0; // @[DCache.scala 126:50]
      end
    end else if (update & updateway1) begin // @[DCache.scala 127:36]
      if (5'h12 == index_addr) begin // @[DCache.scala 127:52]
        d1_18 <= 1'h0; // @[DCache.scala 127:52]
      end
    end else if (way1write) begin // @[DCache.scala 128:25]
      d1_18 <= 5'h12 == index_addr | d1_18;
    end
    if (reset) begin // @[DCache.scala 53:26]
      d1_19 <= 1'h0; // @[DCache.scala 53:26]
    end else if (state == 3'h4) begin // @[DCache.scala 126:35]
      if (5'h13 == fence_cnt) begin // @[DCache.scala 126:50]
        d1_19 <= 1'h0; // @[DCache.scala 126:50]
      end
    end else if (update & updateway1) begin // @[DCache.scala 127:36]
      if (5'h13 == index_addr) begin // @[DCache.scala 127:52]
        d1_19 <= 1'h0; // @[DCache.scala 127:52]
      end
    end else if (way1write) begin // @[DCache.scala 128:25]
      d1_19 <= 5'h13 == index_addr | d1_19;
    end
    if (reset) begin // @[DCache.scala 53:26]
      d1_20 <= 1'h0; // @[DCache.scala 53:26]
    end else if (state == 3'h4) begin // @[DCache.scala 126:35]
      if (5'h14 == fence_cnt) begin // @[DCache.scala 126:50]
        d1_20 <= 1'h0; // @[DCache.scala 126:50]
      end
    end else if (update & updateway1) begin // @[DCache.scala 127:36]
      if (5'h14 == index_addr) begin // @[DCache.scala 127:52]
        d1_20 <= 1'h0; // @[DCache.scala 127:52]
      end
    end else if (way1write) begin // @[DCache.scala 128:25]
      d1_20 <= 5'h14 == index_addr | d1_20;
    end
    if (reset) begin // @[DCache.scala 53:26]
      d1_21 <= 1'h0; // @[DCache.scala 53:26]
    end else if (state == 3'h4) begin // @[DCache.scala 126:35]
      if (5'h15 == fence_cnt) begin // @[DCache.scala 126:50]
        d1_21 <= 1'h0; // @[DCache.scala 126:50]
      end
    end else if (update & updateway1) begin // @[DCache.scala 127:36]
      if (5'h15 == index_addr) begin // @[DCache.scala 127:52]
        d1_21 <= 1'h0; // @[DCache.scala 127:52]
      end
    end else if (way1write) begin // @[DCache.scala 128:25]
      d1_21 <= 5'h15 == index_addr | d1_21;
    end
    if (reset) begin // @[DCache.scala 53:26]
      d1_22 <= 1'h0; // @[DCache.scala 53:26]
    end else if (state == 3'h4) begin // @[DCache.scala 126:35]
      if (5'h16 == fence_cnt) begin // @[DCache.scala 126:50]
        d1_22 <= 1'h0; // @[DCache.scala 126:50]
      end
    end else if (update & updateway1) begin // @[DCache.scala 127:36]
      if (5'h16 == index_addr) begin // @[DCache.scala 127:52]
        d1_22 <= 1'h0; // @[DCache.scala 127:52]
      end
    end else if (way1write) begin // @[DCache.scala 128:25]
      d1_22 <= 5'h16 == index_addr | d1_22;
    end
    if (reset) begin // @[DCache.scala 53:26]
      d1_23 <= 1'h0; // @[DCache.scala 53:26]
    end else if (state == 3'h4) begin // @[DCache.scala 126:35]
      if (5'h17 == fence_cnt) begin // @[DCache.scala 126:50]
        d1_23 <= 1'h0; // @[DCache.scala 126:50]
      end
    end else if (update & updateway1) begin // @[DCache.scala 127:36]
      if (5'h17 == index_addr) begin // @[DCache.scala 127:52]
        d1_23 <= 1'h0; // @[DCache.scala 127:52]
      end
    end else if (way1write) begin // @[DCache.scala 128:25]
      d1_23 <= 5'h17 == index_addr | d1_23;
    end
    if (reset) begin // @[DCache.scala 53:26]
      d1_24 <= 1'h0; // @[DCache.scala 53:26]
    end else if (state == 3'h4) begin // @[DCache.scala 126:35]
      if (5'h18 == fence_cnt) begin // @[DCache.scala 126:50]
        d1_24 <= 1'h0; // @[DCache.scala 126:50]
      end
    end else if (update & updateway1) begin // @[DCache.scala 127:36]
      if (5'h18 == index_addr) begin // @[DCache.scala 127:52]
        d1_24 <= 1'h0; // @[DCache.scala 127:52]
      end
    end else if (way1write) begin // @[DCache.scala 128:25]
      d1_24 <= 5'h18 == index_addr | d1_24;
    end
    if (reset) begin // @[DCache.scala 53:26]
      d1_25 <= 1'h0; // @[DCache.scala 53:26]
    end else if (state == 3'h4) begin // @[DCache.scala 126:35]
      if (5'h19 == fence_cnt) begin // @[DCache.scala 126:50]
        d1_25 <= 1'h0; // @[DCache.scala 126:50]
      end
    end else if (update & updateway1) begin // @[DCache.scala 127:36]
      if (5'h19 == index_addr) begin // @[DCache.scala 127:52]
        d1_25 <= 1'h0; // @[DCache.scala 127:52]
      end
    end else if (way1write) begin // @[DCache.scala 128:25]
      d1_25 <= 5'h19 == index_addr | d1_25;
    end
    if (reset) begin // @[DCache.scala 53:26]
      d1_26 <= 1'h0; // @[DCache.scala 53:26]
    end else if (state == 3'h4) begin // @[DCache.scala 126:35]
      if (5'h1a == fence_cnt) begin // @[DCache.scala 126:50]
        d1_26 <= 1'h0; // @[DCache.scala 126:50]
      end
    end else if (update & updateway1) begin // @[DCache.scala 127:36]
      if (5'h1a == index_addr) begin // @[DCache.scala 127:52]
        d1_26 <= 1'h0; // @[DCache.scala 127:52]
      end
    end else if (way1write) begin // @[DCache.scala 128:25]
      d1_26 <= 5'h1a == index_addr | d1_26;
    end
    if (reset) begin // @[DCache.scala 53:26]
      d1_27 <= 1'h0; // @[DCache.scala 53:26]
    end else if (state == 3'h4) begin // @[DCache.scala 126:35]
      if (5'h1b == fence_cnt) begin // @[DCache.scala 126:50]
        d1_27 <= 1'h0; // @[DCache.scala 126:50]
      end
    end else if (update & updateway1) begin // @[DCache.scala 127:36]
      if (5'h1b == index_addr) begin // @[DCache.scala 127:52]
        d1_27 <= 1'h0; // @[DCache.scala 127:52]
      end
    end else if (way1write) begin // @[DCache.scala 128:25]
      d1_27 <= 5'h1b == index_addr | d1_27;
    end
    if (reset) begin // @[DCache.scala 53:26]
      d1_28 <= 1'h0; // @[DCache.scala 53:26]
    end else if (state == 3'h4) begin // @[DCache.scala 126:35]
      if (5'h1c == fence_cnt) begin // @[DCache.scala 126:50]
        d1_28 <= 1'h0; // @[DCache.scala 126:50]
      end
    end else if (update & updateway1) begin // @[DCache.scala 127:36]
      if (5'h1c == index_addr) begin // @[DCache.scala 127:52]
        d1_28 <= 1'h0; // @[DCache.scala 127:52]
      end
    end else if (way1write) begin // @[DCache.scala 128:25]
      d1_28 <= 5'h1c == index_addr | d1_28;
    end
    if (reset) begin // @[DCache.scala 53:26]
      d1_29 <= 1'h0; // @[DCache.scala 53:26]
    end else if (state == 3'h4) begin // @[DCache.scala 126:35]
      if (5'h1d == fence_cnt) begin // @[DCache.scala 126:50]
        d1_29 <= 1'h0; // @[DCache.scala 126:50]
      end
    end else if (update & updateway1) begin // @[DCache.scala 127:36]
      if (5'h1d == index_addr) begin // @[DCache.scala 127:52]
        d1_29 <= 1'h0; // @[DCache.scala 127:52]
      end
    end else if (way1write) begin // @[DCache.scala 128:25]
      d1_29 <= 5'h1d == index_addr | d1_29;
    end
    if (reset) begin // @[DCache.scala 53:26]
      d1_30 <= 1'h0; // @[DCache.scala 53:26]
    end else if (state == 3'h4) begin // @[DCache.scala 126:35]
      if (5'h1e == fence_cnt) begin // @[DCache.scala 126:50]
        d1_30 <= 1'h0; // @[DCache.scala 126:50]
      end
    end else if (update & updateway1) begin // @[DCache.scala 127:36]
      if (5'h1e == index_addr) begin // @[DCache.scala 127:52]
        d1_30 <= 1'h0; // @[DCache.scala 127:52]
      end
    end else if (way1write) begin // @[DCache.scala 128:25]
      d1_30 <= 5'h1e == index_addr | d1_30;
    end
    if (reset) begin // @[DCache.scala 53:26]
      d1_31 <= 1'h0; // @[DCache.scala 53:26]
    end else if (state == 3'h4) begin // @[DCache.scala 126:35]
      if (5'h1f == fence_cnt) begin // @[DCache.scala 126:50]
        d1_31 <= 1'h0; // @[DCache.scala 126:50]
      end
    end else if (update & updateway1) begin // @[DCache.scala 127:36]
      if (5'h1f == index_addr) begin // @[DCache.scala 127:52]
        d1_31 <= 1'h0; // @[DCache.scala 127:52]
      end
    end else if (way1write) begin // @[DCache.scala 128:25]
      d1_31 <= 5'h1f == index_addr | d1_31;
    end
    if (reset) begin // @[DCache.scala 54:26]
      age1_0 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h0 == index_addr) begin // @[DCache.scala 81:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 81:28]
        age1_0 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 81:28]
        age1_0 <= age1_31; // @[DCache.scala 81:28]
      end else begin
        age1_0 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 54:26]
      age1_1 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h1 == index_addr) begin // @[DCache.scala 81:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 81:28]
        age1_1 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 81:28]
        age1_1 <= age1_31; // @[DCache.scala 81:28]
      end else begin
        age1_1 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 54:26]
      age1_2 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h2 == index_addr) begin // @[DCache.scala 81:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 81:28]
        age1_2 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 81:28]
        age1_2 <= age1_31; // @[DCache.scala 81:28]
      end else begin
        age1_2 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 54:26]
      age1_3 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h3 == index_addr) begin // @[DCache.scala 81:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 81:28]
        age1_3 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 81:28]
        age1_3 <= age1_31; // @[DCache.scala 81:28]
      end else begin
        age1_3 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 54:26]
      age1_4 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h4 == index_addr) begin // @[DCache.scala 81:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 81:28]
        age1_4 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 81:28]
        age1_4 <= age1_31; // @[DCache.scala 81:28]
      end else begin
        age1_4 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 54:26]
      age1_5 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h5 == index_addr) begin // @[DCache.scala 81:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 81:28]
        age1_5 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 81:28]
        age1_5 <= age1_31; // @[DCache.scala 81:28]
      end else begin
        age1_5 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 54:26]
      age1_6 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h6 == index_addr) begin // @[DCache.scala 81:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 81:28]
        age1_6 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 81:28]
        age1_6 <= age1_31; // @[DCache.scala 81:28]
      end else begin
        age1_6 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 54:26]
      age1_7 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h7 == index_addr) begin // @[DCache.scala 81:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 81:28]
        age1_7 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 81:28]
        age1_7 <= age1_31; // @[DCache.scala 81:28]
      end else begin
        age1_7 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 54:26]
      age1_8 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h8 == index_addr) begin // @[DCache.scala 81:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 81:28]
        age1_8 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 81:28]
        age1_8 <= age1_31; // @[DCache.scala 81:28]
      end else begin
        age1_8 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 54:26]
      age1_9 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h9 == index_addr) begin // @[DCache.scala 81:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 81:28]
        age1_9 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 81:28]
        age1_9 <= age1_31; // @[DCache.scala 81:28]
      end else begin
        age1_9 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 54:26]
      age1_10 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'ha == index_addr) begin // @[DCache.scala 81:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 81:28]
        age1_10 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 81:28]
        age1_10 <= age1_31; // @[DCache.scala 81:28]
      end else begin
        age1_10 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 54:26]
      age1_11 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'hb == index_addr) begin // @[DCache.scala 81:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 81:28]
        age1_11 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 81:28]
        age1_11 <= age1_31; // @[DCache.scala 81:28]
      end else begin
        age1_11 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 54:26]
      age1_12 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'hc == index_addr) begin // @[DCache.scala 81:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 81:28]
        age1_12 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 81:28]
        age1_12 <= age1_31; // @[DCache.scala 81:28]
      end else begin
        age1_12 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 54:26]
      age1_13 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'hd == index_addr) begin // @[DCache.scala 81:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 81:28]
        age1_13 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 81:28]
        age1_13 <= age1_31; // @[DCache.scala 81:28]
      end else begin
        age1_13 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 54:26]
      age1_14 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'he == index_addr) begin // @[DCache.scala 81:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 81:28]
        age1_14 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 81:28]
        age1_14 <= age1_31; // @[DCache.scala 81:28]
      end else begin
        age1_14 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 54:26]
      age1_15 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'hf == index_addr) begin // @[DCache.scala 81:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 81:28]
        age1_15 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 81:28]
        age1_15 <= age1_31; // @[DCache.scala 81:28]
      end else begin
        age1_15 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 54:26]
      age1_16 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h10 == index_addr) begin // @[DCache.scala 81:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 81:28]
        age1_16 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 81:28]
        age1_16 <= age1_31; // @[DCache.scala 81:28]
      end else begin
        age1_16 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 54:26]
      age1_17 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h11 == index_addr) begin // @[DCache.scala 81:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 81:28]
        age1_17 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 81:28]
        age1_17 <= age1_31; // @[DCache.scala 81:28]
      end else begin
        age1_17 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 54:26]
      age1_18 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h12 == index_addr) begin // @[DCache.scala 81:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 81:28]
        age1_18 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 81:28]
        age1_18 <= age1_31; // @[DCache.scala 81:28]
      end else begin
        age1_18 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 54:26]
      age1_19 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h13 == index_addr) begin // @[DCache.scala 81:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 81:28]
        age1_19 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 81:28]
        age1_19 <= age1_31; // @[DCache.scala 81:28]
      end else begin
        age1_19 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 54:26]
      age1_20 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h14 == index_addr) begin // @[DCache.scala 81:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 81:28]
        age1_20 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 81:28]
        age1_20 <= age1_31; // @[DCache.scala 81:28]
      end else begin
        age1_20 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 54:26]
      age1_21 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h15 == index_addr) begin // @[DCache.scala 81:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 81:28]
        age1_21 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 81:28]
        age1_21 <= age1_31; // @[DCache.scala 81:28]
      end else begin
        age1_21 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 54:26]
      age1_22 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h16 == index_addr) begin // @[DCache.scala 81:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 81:28]
        age1_22 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 81:28]
        age1_22 <= age1_31; // @[DCache.scala 81:28]
      end else begin
        age1_22 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 54:26]
      age1_23 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h17 == index_addr) begin // @[DCache.scala 81:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 81:28]
        age1_23 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 81:28]
        age1_23 <= age1_31; // @[DCache.scala 81:28]
      end else begin
        age1_23 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 54:26]
      age1_24 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h18 == index_addr) begin // @[DCache.scala 81:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 81:28]
        age1_24 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 81:28]
        age1_24 <= age1_31; // @[DCache.scala 81:28]
      end else begin
        age1_24 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 54:26]
      age1_25 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h19 == index_addr) begin // @[DCache.scala 81:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 81:28]
        age1_25 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 81:28]
        age1_25 <= age1_31; // @[DCache.scala 81:28]
      end else begin
        age1_25 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 54:26]
      age1_26 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h1a == index_addr) begin // @[DCache.scala 81:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 81:28]
        age1_26 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 81:28]
        age1_26 <= age1_31; // @[DCache.scala 81:28]
      end else begin
        age1_26 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 54:26]
      age1_27 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h1b == index_addr) begin // @[DCache.scala 81:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 81:28]
        age1_27 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 81:28]
        age1_27 <= age1_31; // @[DCache.scala 81:28]
      end else begin
        age1_27 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 54:26]
      age1_28 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h1c == index_addr) begin // @[DCache.scala 81:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 81:28]
        age1_28 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 81:28]
        age1_28 <= age1_31; // @[DCache.scala 81:28]
      end else begin
        age1_28 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 54:26]
      age1_29 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h1d == index_addr) begin // @[DCache.scala 81:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 81:28]
        age1_29 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 81:28]
        age1_29 <= age1_31; // @[DCache.scala 81:28]
      end else begin
        age1_29 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 54:26]
      age1_30 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h1e == index_addr) begin // @[DCache.scala 81:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 81:28]
        age1_30 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 81:28]
        age1_30 <= age1_31; // @[DCache.scala 81:28]
      end else begin
        age1_30 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 54:26]
      age1_31 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h1f == index_addr) begin // @[DCache.scala 81:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 81:28]
        age1_31 <= hit1;
      end else if (!(5'h1f == index_addr)) begin // @[DCache.scala 81:28]
        age1_31 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      tag1_0 <= 53'h0; // @[DCache.scala 55:26]
    end else if (5'h0 == index_addr) begin // @[DCache.scala 144:26]
      if (_T_20) begin // @[DCache.scala 144:32]
        tag1_0 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 63:28]
        tag1_0 <= tag1_31; // @[DCache.scala 63:28]
      end else begin
        tag1_0 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      tag1_1 <= 53'h0; // @[DCache.scala 55:26]
    end else if (5'h1 == index_addr) begin // @[DCache.scala 144:26]
      if (_T_20) begin // @[DCache.scala 144:32]
        tag1_1 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 63:28]
        tag1_1 <= tag1_31; // @[DCache.scala 63:28]
      end else begin
        tag1_1 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      tag1_2 <= 53'h0; // @[DCache.scala 55:26]
    end else if (5'h2 == index_addr) begin // @[DCache.scala 144:26]
      if (_T_20) begin // @[DCache.scala 144:32]
        tag1_2 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 63:28]
        tag1_2 <= tag1_31; // @[DCache.scala 63:28]
      end else begin
        tag1_2 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      tag1_3 <= 53'h0; // @[DCache.scala 55:26]
    end else if (5'h3 == index_addr) begin // @[DCache.scala 144:26]
      if (_T_20) begin // @[DCache.scala 144:32]
        tag1_3 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 63:28]
        tag1_3 <= tag1_31; // @[DCache.scala 63:28]
      end else begin
        tag1_3 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      tag1_4 <= 53'h0; // @[DCache.scala 55:26]
    end else if (5'h4 == index_addr) begin // @[DCache.scala 144:26]
      if (_T_20) begin // @[DCache.scala 144:32]
        tag1_4 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 63:28]
        tag1_4 <= tag1_31; // @[DCache.scala 63:28]
      end else begin
        tag1_4 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      tag1_5 <= 53'h0; // @[DCache.scala 55:26]
    end else if (5'h5 == index_addr) begin // @[DCache.scala 144:26]
      if (_T_20) begin // @[DCache.scala 144:32]
        tag1_5 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 63:28]
        tag1_5 <= tag1_31; // @[DCache.scala 63:28]
      end else begin
        tag1_5 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      tag1_6 <= 53'h0; // @[DCache.scala 55:26]
    end else if (5'h6 == index_addr) begin // @[DCache.scala 144:26]
      if (_T_20) begin // @[DCache.scala 144:32]
        tag1_6 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 63:28]
        tag1_6 <= tag1_31; // @[DCache.scala 63:28]
      end else begin
        tag1_6 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      tag1_7 <= 53'h0; // @[DCache.scala 55:26]
    end else if (5'h7 == index_addr) begin // @[DCache.scala 144:26]
      if (_T_20) begin // @[DCache.scala 144:32]
        tag1_7 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 63:28]
        tag1_7 <= tag1_31; // @[DCache.scala 63:28]
      end else begin
        tag1_7 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      tag1_8 <= 53'h0; // @[DCache.scala 55:26]
    end else if (5'h8 == index_addr) begin // @[DCache.scala 144:26]
      if (_T_20) begin // @[DCache.scala 144:32]
        tag1_8 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 63:28]
        tag1_8 <= tag1_31; // @[DCache.scala 63:28]
      end else begin
        tag1_8 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      tag1_9 <= 53'h0; // @[DCache.scala 55:26]
    end else if (5'h9 == index_addr) begin // @[DCache.scala 144:26]
      if (_T_20) begin // @[DCache.scala 144:32]
        tag1_9 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 63:28]
        tag1_9 <= tag1_31; // @[DCache.scala 63:28]
      end else begin
        tag1_9 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      tag1_10 <= 53'h0; // @[DCache.scala 55:26]
    end else if (5'ha == index_addr) begin // @[DCache.scala 144:26]
      if (_T_20) begin // @[DCache.scala 144:32]
        tag1_10 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 63:28]
        tag1_10 <= tag1_31; // @[DCache.scala 63:28]
      end else begin
        tag1_10 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      tag1_11 <= 53'h0; // @[DCache.scala 55:26]
    end else if (5'hb == index_addr) begin // @[DCache.scala 144:26]
      if (_T_20) begin // @[DCache.scala 144:32]
        tag1_11 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 63:28]
        tag1_11 <= tag1_31; // @[DCache.scala 63:28]
      end else begin
        tag1_11 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      tag1_12 <= 53'h0; // @[DCache.scala 55:26]
    end else if (5'hc == index_addr) begin // @[DCache.scala 144:26]
      if (_T_20) begin // @[DCache.scala 144:32]
        tag1_12 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 63:28]
        tag1_12 <= tag1_31; // @[DCache.scala 63:28]
      end else begin
        tag1_12 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      tag1_13 <= 53'h0; // @[DCache.scala 55:26]
    end else if (5'hd == index_addr) begin // @[DCache.scala 144:26]
      if (_T_20) begin // @[DCache.scala 144:32]
        tag1_13 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 63:28]
        tag1_13 <= tag1_31; // @[DCache.scala 63:28]
      end else begin
        tag1_13 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      tag1_14 <= 53'h0; // @[DCache.scala 55:26]
    end else if (5'he == index_addr) begin // @[DCache.scala 144:26]
      if (_T_20) begin // @[DCache.scala 144:32]
        tag1_14 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 63:28]
        tag1_14 <= tag1_31; // @[DCache.scala 63:28]
      end else begin
        tag1_14 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      tag1_15 <= 53'h0; // @[DCache.scala 55:26]
    end else if (5'hf == index_addr) begin // @[DCache.scala 144:26]
      if (_T_20) begin // @[DCache.scala 144:32]
        tag1_15 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 63:28]
        tag1_15 <= tag1_31; // @[DCache.scala 63:28]
      end else begin
        tag1_15 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      tag1_16 <= 53'h0; // @[DCache.scala 55:26]
    end else if (5'h10 == index_addr) begin // @[DCache.scala 144:26]
      if (_T_20) begin // @[DCache.scala 144:32]
        tag1_16 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 63:28]
        tag1_16 <= tag1_31; // @[DCache.scala 63:28]
      end else begin
        tag1_16 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      tag1_17 <= 53'h0; // @[DCache.scala 55:26]
    end else if (5'h11 == index_addr) begin // @[DCache.scala 144:26]
      if (_T_20) begin // @[DCache.scala 144:32]
        tag1_17 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 63:28]
        tag1_17 <= tag1_31; // @[DCache.scala 63:28]
      end else begin
        tag1_17 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      tag1_18 <= 53'h0; // @[DCache.scala 55:26]
    end else if (5'h12 == index_addr) begin // @[DCache.scala 144:26]
      if (_T_20) begin // @[DCache.scala 144:32]
        tag1_18 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 63:28]
        tag1_18 <= tag1_31; // @[DCache.scala 63:28]
      end else begin
        tag1_18 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      tag1_19 <= 53'h0; // @[DCache.scala 55:26]
    end else if (5'h13 == index_addr) begin // @[DCache.scala 144:26]
      if (_T_20) begin // @[DCache.scala 144:32]
        tag1_19 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 63:28]
        tag1_19 <= tag1_31; // @[DCache.scala 63:28]
      end else begin
        tag1_19 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      tag1_20 <= 53'h0; // @[DCache.scala 55:26]
    end else if (5'h14 == index_addr) begin // @[DCache.scala 144:26]
      if (_T_20) begin // @[DCache.scala 144:32]
        tag1_20 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 63:28]
        tag1_20 <= tag1_31; // @[DCache.scala 63:28]
      end else begin
        tag1_20 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      tag1_21 <= 53'h0; // @[DCache.scala 55:26]
    end else if (5'h15 == index_addr) begin // @[DCache.scala 144:26]
      if (_T_20) begin // @[DCache.scala 144:32]
        tag1_21 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 63:28]
        tag1_21 <= tag1_31; // @[DCache.scala 63:28]
      end else begin
        tag1_21 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      tag1_22 <= 53'h0; // @[DCache.scala 55:26]
    end else if (5'h16 == index_addr) begin // @[DCache.scala 144:26]
      if (_T_20) begin // @[DCache.scala 144:32]
        tag1_22 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 63:28]
        tag1_22 <= tag1_31; // @[DCache.scala 63:28]
      end else begin
        tag1_22 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      tag1_23 <= 53'h0; // @[DCache.scala 55:26]
    end else if (5'h17 == index_addr) begin // @[DCache.scala 144:26]
      if (_T_20) begin // @[DCache.scala 144:32]
        tag1_23 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 63:28]
        tag1_23 <= tag1_31; // @[DCache.scala 63:28]
      end else begin
        tag1_23 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      tag1_24 <= 53'h0; // @[DCache.scala 55:26]
    end else if (5'h18 == index_addr) begin // @[DCache.scala 144:26]
      if (_T_20) begin // @[DCache.scala 144:32]
        tag1_24 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 63:28]
        tag1_24 <= tag1_31; // @[DCache.scala 63:28]
      end else begin
        tag1_24 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      tag1_25 <= 53'h0; // @[DCache.scala 55:26]
    end else if (5'h19 == index_addr) begin // @[DCache.scala 144:26]
      if (_T_20) begin // @[DCache.scala 144:32]
        tag1_25 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 63:28]
        tag1_25 <= tag1_31; // @[DCache.scala 63:28]
      end else begin
        tag1_25 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      tag1_26 <= 53'h0; // @[DCache.scala 55:26]
    end else if (5'h1a == index_addr) begin // @[DCache.scala 144:26]
      if (_T_20) begin // @[DCache.scala 144:32]
        tag1_26 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 63:28]
        tag1_26 <= tag1_31; // @[DCache.scala 63:28]
      end else begin
        tag1_26 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      tag1_27 <= 53'h0; // @[DCache.scala 55:26]
    end else if (5'h1b == index_addr) begin // @[DCache.scala 144:26]
      if (_T_20) begin // @[DCache.scala 144:32]
        tag1_27 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 63:28]
        tag1_27 <= tag1_31; // @[DCache.scala 63:28]
      end else begin
        tag1_27 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      tag1_28 <= 53'h0; // @[DCache.scala 55:26]
    end else if (5'h1c == index_addr) begin // @[DCache.scala 144:26]
      if (_T_20) begin // @[DCache.scala 144:32]
        tag1_28 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 63:28]
        tag1_28 <= tag1_31; // @[DCache.scala 63:28]
      end else begin
        tag1_28 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      tag1_29 <= 53'h0; // @[DCache.scala 55:26]
    end else if (5'h1d == index_addr) begin // @[DCache.scala 144:26]
      if (_T_20) begin // @[DCache.scala 144:32]
        tag1_29 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 63:28]
        tag1_29 <= tag1_31; // @[DCache.scala 63:28]
      end else begin
        tag1_29 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      tag1_30 <= 53'h0; // @[DCache.scala 55:26]
    end else if (5'h1e == index_addr) begin // @[DCache.scala 144:26]
      if (_T_20) begin // @[DCache.scala 144:32]
        tag1_30 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 63:28]
        tag1_30 <= tag1_31; // @[DCache.scala 63:28]
      end else begin
        tag1_30 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      tag1_31 <= 53'h0; // @[DCache.scala 55:26]
    end else if (5'h1f == index_addr) begin // @[DCache.scala 144:26]
      if (_T_20) begin // @[DCache.scala 144:32]
        tag1_31 <= tag_addr;
      end else if (!(5'h1f == index_addr)) begin // @[DCache.scala 63:28]
        tag1_31 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      block1_0 <= 512'h0; // @[DCache.scala 56:26]
    end else if (5'h0 == index_addr) begin // @[DCache.scala 143:26]
      if (_T_20) begin // @[DCache.scala 143:32]
        block1_0 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 143:72]
        block1_0 <= block1_after_write;
      end else begin
        block1_0 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      block1_1 <= 512'h0; // @[DCache.scala 56:26]
    end else if (5'h1 == index_addr) begin // @[DCache.scala 143:26]
      if (_T_20) begin // @[DCache.scala 143:32]
        block1_1 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 143:72]
        block1_1 <= block1_after_write;
      end else begin
        block1_1 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      block1_2 <= 512'h0; // @[DCache.scala 56:26]
    end else if (5'h2 == index_addr) begin // @[DCache.scala 143:26]
      if (_T_20) begin // @[DCache.scala 143:32]
        block1_2 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 143:72]
        block1_2 <= block1_after_write;
      end else begin
        block1_2 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      block1_3 <= 512'h0; // @[DCache.scala 56:26]
    end else if (5'h3 == index_addr) begin // @[DCache.scala 143:26]
      if (_T_20) begin // @[DCache.scala 143:32]
        block1_3 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 143:72]
        block1_3 <= block1_after_write;
      end else begin
        block1_3 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      block1_4 <= 512'h0; // @[DCache.scala 56:26]
    end else if (5'h4 == index_addr) begin // @[DCache.scala 143:26]
      if (_T_20) begin // @[DCache.scala 143:32]
        block1_4 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 143:72]
        block1_4 <= block1_after_write;
      end else begin
        block1_4 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      block1_5 <= 512'h0; // @[DCache.scala 56:26]
    end else if (5'h5 == index_addr) begin // @[DCache.scala 143:26]
      if (_T_20) begin // @[DCache.scala 143:32]
        block1_5 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 143:72]
        block1_5 <= block1_after_write;
      end else begin
        block1_5 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      block1_6 <= 512'h0; // @[DCache.scala 56:26]
    end else if (5'h6 == index_addr) begin // @[DCache.scala 143:26]
      if (_T_20) begin // @[DCache.scala 143:32]
        block1_6 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 143:72]
        block1_6 <= block1_after_write;
      end else begin
        block1_6 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      block1_7 <= 512'h0; // @[DCache.scala 56:26]
    end else if (5'h7 == index_addr) begin // @[DCache.scala 143:26]
      if (_T_20) begin // @[DCache.scala 143:32]
        block1_7 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 143:72]
        block1_7 <= block1_after_write;
      end else begin
        block1_7 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      block1_8 <= 512'h0; // @[DCache.scala 56:26]
    end else if (5'h8 == index_addr) begin // @[DCache.scala 143:26]
      if (_T_20) begin // @[DCache.scala 143:32]
        block1_8 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 143:72]
        block1_8 <= block1_after_write;
      end else begin
        block1_8 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      block1_9 <= 512'h0; // @[DCache.scala 56:26]
    end else if (5'h9 == index_addr) begin // @[DCache.scala 143:26]
      if (_T_20) begin // @[DCache.scala 143:32]
        block1_9 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 143:72]
        block1_9 <= block1_after_write;
      end else begin
        block1_9 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      block1_10 <= 512'h0; // @[DCache.scala 56:26]
    end else if (5'ha == index_addr) begin // @[DCache.scala 143:26]
      if (_T_20) begin // @[DCache.scala 143:32]
        block1_10 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 143:72]
        block1_10 <= block1_after_write;
      end else begin
        block1_10 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      block1_11 <= 512'h0; // @[DCache.scala 56:26]
    end else if (5'hb == index_addr) begin // @[DCache.scala 143:26]
      if (_T_20) begin // @[DCache.scala 143:32]
        block1_11 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 143:72]
        block1_11 <= block1_after_write;
      end else begin
        block1_11 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      block1_12 <= 512'h0; // @[DCache.scala 56:26]
    end else if (5'hc == index_addr) begin // @[DCache.scala 143:26]
      if (_T_20) begin // @[DCache.scala 143:32]
        block1_12 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 143:72]
        block1_12 <= block1_after_write;
      end else begin
        block1_12 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      block1_13 <= 512'h0; // @[DCache.scala 56:26]
    end else if (5'hd == index_addr) begin // @[DCache.scala 143:26]
      if (_T_20) begin // @[DCache.scala 143:32]
        block1_13 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 143:72]
        block1_13 <= block1_after_write;
      end else begin
        block1_13 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      block1_14 <= 512'h0; // @[DCache.scala 56:26]
    end else if (5'he == index_addr) begin // @[DCache.scala 143:26]
      if (_T_20) begin // @[DCache.scala 143:32]
        block1_14 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 143:72]
        block1_14 <= block1_after_write;
      end else begin
        block1_14 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      block1_15 <= 512'h0; // @[DCache.scala 56:26]
    end else if (5'hf == index_addr) begin // @[DCache.scala 143:26]
      if (_T_20) begin // @[DCache.scala 143:32]
        block1_15 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 143:72]
        block1_15 <= block1_after_write;
      end else begin
        block1_15 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      block1_16 <= 512'h0; // @[DCache.scala 56:26]
    end else if (5'h10 == index_addr) begin // @[DCache.scala 143:26]
      if (_T_20) begin // @[DCache.scala 143:32]
        block1_16 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 143:72]
        block1_16 <= block1_after_write;
      end else begin
        block1_16 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      block1_17 <= 512'h0; // @[DCache.scala 56:26]
    end else if (5'h11 == index_addr) begin // @[DCache.scala 143:26]
      if (_T_20) begin // @[DCache.scala 143:32]
        block1_17 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 143:72]
        block1_17 <= block1_after_write;
      end else begin
        block1_17 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      block1_18 <= 512'h0; // @[DCache.scala 56:26]
    end else if (5'h12 == index_addr) begin // @[DCache.scala 143:26]
      if (_T_20) begin // @[DCache.scala 143:32]
        block1_18 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 143:72]
        block1_18 <= block1_after_write;
      end else begin
        block1_18 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      block1_19 <= 512'h0; // @[DCache.scala 56:26]
    end else if (5'h13 == index_addr) begin // @[DCache.scala 143:26]
      if (_T_20) begin // @[DCache.scala 143:32]
        block1_19 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 143:72]
        block1_19 <= block1_after_write;
      end else begin
        block1_19 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      block1_20 <= 512'h0; // @[DCache.scala 56:26]
    end else if (5'h14 == index_addr) begin // @[DCache.scala 143:26]
      if (_T_20) begin // @[DCache.scala 143:32]
        block1_20 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 143:72]
        block1_20 <= block1_after_write;
      end else begin
        block1_20 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      block1_21 <= 512'h0; // @[DCache.scala 56:26]
    end else if (5'h15 == index_addr) begin // @[DCache.scala 143:26]
      if (_T_20) begin // @[DCache.scala 143:32]
        block1_21 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 143:72]
        block1_21 <= block1_after_write;
      end else begin
        block1_21 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      block1_22 <= 512'h0; // @[DCache.scala 56:26]
    end else if (5'h16 == index_addr) begin // @[DCache.scala 143:26]
      if (_T_20) begin // @[DCache.scala 143:32]
        block1_22 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 143:72]
        block1_22 <= block1_after_write;
      end else begin
        block1_22 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      block1_23 <= 512'h0; // @[DCache.scala 56:26]
    end else if (5'h17 == index_addr) begin // @[DCache.scala 143:26]
      if (_T_20) begin // @[DCache.scala 143:32]
        block1_23 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 143:72]
        block1_23 <= block1_after_write;
      end else begin
        block1_23 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      block1_24 <= 512'h0; // @[DCache.scala 56:26]
    end else if (5'h18 == index_addr) begin // @[DCache.scala 143:26]
      if (_T_20) begin // @[DCache.scala 143:32]
        block1_24 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 143:72]
        block1_24 <= block1_after_write;
      end else begin
        block1_24 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      block1_25 <= 512'h0; // @[DCache.scala 56:26]
    end else if (5'h19 == index_addr) begin // @[DCache.scala 143:26]
      if (_T_20) begin // @[DCache.scala 143:32]
        block1_25 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 143:72]
        block1_25 <= block1_after_write;
      end else begin
        block1_25 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      block1_26 <= 512'h0; // @[DCache.scala 56:26]
    end else if (5'h1a == index_addr) begin // @[DCache.scala 143:26]
      if (_T_20) begin // @[DCache.scala 143:32]
        block1_26 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 143:72]
        block1_26 <= block1_after_write;
      end else begin
        block1_26 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      block1_27 <= 512'h0; // @[DCache.scala 56:26]
    end else if (5'h1b == index_addr) begin // @[DCache.scala 143:26]
      if (_T_20) begin // @[DCache.scala 143:32]
        block1_27 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 143:72]
        block1_27 <= block1_after_write;
      end else begin
        block1_27 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      block1_28 <= 512'h0; // @[DCache.scala 56:26]
    end else if (5'h1c == index_addr) begin // @[DCache.scala 143:26]
      if (_T_20) begin // @[DCache.scala 143:32]
        block1_28 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 143:72]
        block1_28 <= block1_after_write;
      end else begin
        block1_28 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      block1_29 <= 512'h0; // @[DCache.scala 56:26]
    end else if (5'h1d == index_addr) begin // @[DCache.scala 143:26]
      if (_T_20) begin // @[DCache.scala 143:32]
        block1_29 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 143:72]
        block1_29 <= block1_after_write;
      end else begin
        block1_29 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      block1_30 <= 512'h0; // @[DCache.scala 56:26]
    end else if (5'h1e == index_addr) begin // @[DCache.scala 143:26]
      if (_T_20) begin // @[DCache.scala 143:32]
        block1_30 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 143:72]
        block1_30 <= block1_after_write;
      end else begin
        block1_30 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      block1_31 <= 512'h0; // @[DCache.scala 56:26]
    end else if (5'h1f == index_addr) begin // @[DCache.scala 143:26]
      if (_T_20) begin // @[DCache.scala 143:32]
        block1_31 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 143:72]
        block1_31 <= block1_after_write;
      end else begin
        block1_31 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 57:26]
      v2_0 <= 1'h0; // @[DCache.scala 57:26]
    end else if (5'h0 == index_addr) begin // @[DCache.scala 148:26]
      v2_0 <= _T_22 | _GEN_131; // @[DCache.scala 148:26]
    end
    if (reset) begin // @[DCache.scala 57:26]
      v2_1 <= 1'h0; // @[DCache.scala 57:26]
    end else if (5'h1 == index_addr) begin // @[DCache.scala 148:26]
      v2_1 <= _T_22 | _GEN_131; // @[DCache.scala 148:26]
    end
    if (reset) begin // @[DCache.scala 57:26]
      v2_2 <= 1'h0; // @[DCache.scala 57:26]
    end else if (5'h2 == index_addr) begin // @[DCache.scala 148:26]
      v2_2 <= _T_22 | _GEN_131; // @[DCache.scala 148:26]
    end
    if (reset) begin // @[DCache.scala 57:26]
      v2_3 <= 1'h0; // @[DCache.scala 57:26]
    end else if (5'h3 == index_addr) begin // @[DCache.scala 148:26]
      v2_3 <= _T_22 | _GEN_131; // @[DCache.scala 148:26]
    end
    if (reset) begin // @[DCache.scala 57:26]
      v2_4 <= 1'h0; // @[DCache.scala 57:26]
    end else if (5'h4 == index_addr) begin // @[DCache.scala 148:26]
      v2_4 <= _T_22 | _GEN_131; // @[DCache.scala 148:26]
    end
    if (reset) begin // @[DCache.scala 57:26]
      v2_5 <= 1'h0; // @[DCache.scala 57:26]
    end else if (5'h5 == index_addr) begin // @[DCache.scala 148:26]
      v2_5 <= _T_22 | _GEN_131; // @[DCache.scala 148:26]
    end
    if (reset) begin // @[DCache.scala 57:26]
      v2_6 <= 1'h0; // @[DCache.scala 57:26]
    end else if (5'h6 == index_addr) begin // @[DCache.scala 148:26]
      v2_6 <= _T_22 | _GEN_131; // @[DCache.scala 148:26]
    end
    if (reset) begin // @[DCache.scala 57:26]
      v2_7 <= 1'h0; // @[DCache.scala 57:26]
    end else if (5'h7 == index_addr) begin // @[DCache.scala 148:26]
      v2_7 <= _T_22 | _GEN_131; // @[DCache.scala 148:26]
    end
    if (reset) begin // @[DCache.scala 57:26]
      v2_8 <= 1'h0; // @[DCache.scala 57:26]
    end else if (5'h8 == index_addr) begin // @[DCache.scala 148:26]
      v2_8 <= _T_22 | _GEN_131; // @[DCache.scala 148:26]
    end
    if (reset) begin // @[DCache.scala 57:26]
      v2_9 <= 1'h0; // @[DCache.scala 57:26]
    end else if (5'h9 == index_addr) begin // @[DCache.scala 148:26]
      v2_9 <= _T_22 | _GEN_131; // @[DCache.scala 148:26]
    end
    if (reset) begin // @[DCache.scala 57:26]
      v2_10 <= 1'h0; // @[DCache.scala 57:26]
    end else if (5'ha == index_addr) begin // @[DCache.scala 148:26]
      v2_10 <= _T_22 | _GEN_131; // @[DCache.scala 148:26]
    end
    if (reset) begin // @[DCache.scala 57:26]
      v2_11 <= 1'h0; // @[DCache.scala 57:26]
    end else if (5'hb == index_addr) begin // @[DCache.scala 148:26]
      v2_11 <= _T_22 | _GEN_131; // @[DCache.scala 148:26]
    end
    if (reset) begin // @[DCache.scala 57:26]
      v2_12 <= 1'h0; // @[DCache.scala 57:26]
    end else if (5'hc == index_addr) begin // @[DCache.scala 148:26]
      v2_12 <= _T_22 | _GEN_131; // @[DCache.scala 148:26]
    end
    if (reset) begin // @[DCache.scala 57:26]
      v2_13 <= 1'h0; // @[DCache.scala 57:26]
    end else if (5'hd == index_addr) begin // @[DCache.scala 148:26]
      v2_13 <= _T_22 | _GEN_131; // @[DCache.scala 148:26]
    end
    if (reset) begin // @[DCache.scala 57:26]
      v2_14 <= 1'h0; // @[DCache.scala 57:26]
    end else if (5'he == index_addr) begin // @[DCache.scala 148:26]
      v2_14 <= _T_22 | _GEN_131; // @[DCache.scala 148:26]
    end
    if (reset) begin // @[DCache.scala 57:26]
      v2_15 <= 1'h0; // @[DCache.scala 57:26]
    end else if (5'hf == index_addr) begin // @[DCache.scala 148:26]
      v2_15 <= _T_22 | _GEN_131; // @[DCache.scala 148:26]
    end
    if (reset) begin // @[DCache.scala 57:26]
      v2_16 <= 1'h0; // @[DCache.scala 57:26]
    end else if (5'h10 == index_addr) begin // @[DCache.scala 148:26]
      v2_16 <= _T_22 | _GEN_131; // @[DCache.scala 148:26]
    end
    if (reset) begin // @[DCache.scala 57:26]
      v2_17 <= 1'h0; // @[DCache.scala 57:26]
    end else if (5'h11 == index_addr) begin // @[DCache.scala 148:26]
      v2_17 <= _T_22 | _GEN_131; // @[DCache.scala 148:26]
    end
    if (reset) begin // @[DCache.scala 57:26]
      v2_18 <= 1'h0; // @[DCache.scala 57:26]
    end else if (5'h12 == index_addr) begin // @[DCache.scala 148:26]
      v2_18 <= _T_22 | _GEN_131; // @[DCache.scala 148:26]
    end
    if (reset) begin // @[DCache.scala 57:26]
      v2_19 <= 1'h0; // @[DCache.scala 57:26]
    end else if (5'h13 == index_addr) begin // @[DCache.scala 148:26]
      v2_19 <= _T_22 | _GEN_131; // @[DCache.scala 148:26]
    end
    if (reset) begin // @[DCache.scala 57:26]
      v2_20 <= 1'h0; // @[DCache.scala 57:26]
    end else if (5'h14 == index_addr) begin // @[DCache.scala 148:26]
      v2_20 <= _T_22 | _GEN_131; // @[DCache.scala 148:26]
    end
    if (reset) begin // @[DCache.scala 57:26]
      v2_21 <= 1'h0; // @[DCache.scala 57:26]
    end else if (5'h15 == index_addr) begin // @[DCache.scala 148:26]
      v2_21 <= _T_22 | _GEN_131; // @[DCache.scala 148:26]
    end
    if (reset) begin // @[DCache.scala 57:26]
      v2_22 <= 1'h0; // @[DCache.scala 57:26]
    end else if (5'h16 == index_addr) begin // @[DCache.scala 148:26]
      v2_22 <= _T_22 | _GEN_131; // @[DCache.scala 148:26]
    end
    if (reset) begin // @[DCache.scala 57:26]
      v2_23 <= 1'h0; // @[DCache.scala 57:26]
    end else if (5'h17 == index_addr) begin // @[DCache.scala 148:26]
      v2_23 <= _T_22 | _GEN_131; // @[DCache.scala 148:26]
    end
    if (reset) begin // @[DCache.scala 57:26]
      v2_24 <= 1'h0; // @[DCache.scala 57:26]
    end else if (5'h18 == index_addr) begin // @[DCache.scala 148:26]
      v2_24 <= _T_22 | _GEN_131; // @[DCache.scala 148:26]
    end
    if (reset) begin // @[DCache.scala 57:26]
      v2_25 <= 1'h0; // @[DCache.scala 57:26]
    end else if (5'h19 == index_addr) begin // @[DCache.scala 148:26]
      v2_25 <= _T_22 | _GEN_131; // @[DCache.scala 148:26]
    end
    if (reset) begin // @[DCache.scala 57:26]
      v2_26 <= 1'h0; // @[DCache.scala 57:26]
    end else if (5'h1a == index_addr) begin // @[DCache.scala 148:26]
      v2_26 <= _T_22 | _GEN_131; // @[DCache.scala 148:26]
    end
    if (reset) begin // @[DCache.scala 57:26]
      v2_27 <= 1'h0; // @[DCache.scala 57:26]
    end else if (5'h1b == index_addr) begin // @[DCache.scala 148:26]
      v2_27 <= _T_22 | _GEN_131; // @[DCache.scala 148:26]
    end
    if (reset) begin // @[DCache.scala 57:26]
      v2_28 <= 1'h0; // @[DCache.scala 57:26]
    end else if (5'h1c == index_addr) begin // @[DCache.scala 148:26]
      v2_28 <= _T_22 | _GEN_131; // @[DCache.scala 148:26]
    end
    if (reset) begin // @[DCache.scala 57:26]
      v2_29 <= 1'h0; // @[DCache.scala 57:26]
    end else if (5'h1d == index_addr) begin // @[DCache.scala 148:26]
      v2_29 <= _T_22 | _GEN_131; // @[DCache.scala 148:26]
    end
    if (reset) begin // @[DCache.scala 57:26]
      v2_30 <= 1'h0; // @[DCache.scala 57:26]
    end else if (5'h1e == index_addr) begin // @[DCache.scala 148:26]
      v2_30 <= _T_22 | _GEN_131; // @[DCache.scala 148:26]
    end
    if (reset) begin // @[DCache.scala 57:26]
      v2_31 <= 1'h0; // @[DCache.scala 57:26]
    end else if (5'h1f == index_addr) begin // @[DCache.scala 148:26]
      v2_31 <= _T_22 | _GEN_131; // @[DCache.scala 148:26]
    end
    if (reset) begin // @[DCache.scala 58:26]
      d2_0 <= 1'h0; // @[DCache.scala 58:26]
    end else if (state == 3'h6) begin // @[DCache.scala 130:35]
      if (5'h0 == fence_cnt) begin // @[DCache.scala 130:50]
        d2_0 <= 1'h0; // @[DCache.scala 130:50]
      end
    end else if (update & updateway2) begin // @[DCache.scala 131:36]
      if (5'h0 == index_addr) begin // @[DCache.scala 131:52]
        d2_0 <= 1'h0; // @[DCache.scala 131:52]
      end
    end else if (way2write) begin // @[DCache.scala 132:25]
      d2_0 <= _GEN_1182 | d2_0;
    end
    if (reset) begin // @[DCache.scala 58:26]
      d2_1 <= 1'h0; // @[DCache.scala 58:26]
    end else if (state == 3'h6) begin // @[DCache.scala 130:35]
      if (5'h1 == fence_cnt) begin // @[DCache.scala 130:50]
        d2_1 <= 1'h0; // @[DCache.scala 130:50]
      end
    end else if (update & updateway2) begin // @[DCache.scala 131:36]
      if (5'h1 == index_addr) begin // @[DCache.scala 131:52]
        d2_1 <= 1'h0; // @[DCache.scala 131:52]
      end
    end else if (way2write) begin // @[DCache.scala 132:25]
      d2_1 <= _GEN_1183 | d2_1;
    end
    if (reset) begin // @[DCache.scala 58:26]
      d2_2 <= 1'h0; // @[DCache.scala 58:26]
    end else if (state == 3'h6) begin // @[DCache.scala 130:35]
      if (5'h2 == fence_cnt) begin // @[DCache.scala 130:50]
        d2_2 <= 1'h0; // @[DCache.scala 130:50]
      end
    end else if (update & updateway2) begin // @[DCache.scala 131:36]
      if (5'h2 == index_addr) begin // @[DCache.scala 131:52]
        d2_2 <= 1'h0; // @[DCache.scala 131:52]
      end
    end else if (way2write) begin // @[DCache.scala 132:25]
      d2_2 <= _GEN_1184 | d2_2;
    end
    if (reset) begin // @[DCache.scala 58:26]
      d2_3 <= 1'h0; // @[DCache.scala 58:26]
    end else if (state == 3'h6) begin // @[DCache.scala 130:35]
      if (5'h3 == fence_cnt) begin // @[DCache.scala 130:50]
        d2_3 <= 1'h0; // @[DCache.scala 130:50]
      end
    end else if (update & updateway2) begin // @[DCache.scala 131:36]
      if (5'h3 == index_addr) begin // @[DCache.scala 131:52]
        d2_3 <= 1'h0; // @[DCache.scala 131:52]
      end
    end else if (way2write) begin // @[DCache.scala 132:25]
      d2_3 <= _GEN_1185 | d2_3;
    end
    if (reset) begin // @[DCache.scala 58:26]
      d2_4 <= 1'h0; // @[DCache.scala 58:26]
    end else if (state == 3'h6) begin // @[DCache.scala 130:35]
      if (5'h4 == fence_cnt) begin // @[DCache.scala 130:50]
        d2_4 <= 1'h0; // @[DCache.scala 130:50]
      end
    end else if (update & updateway2) begin // @[DCache.scala 131:36]
      if (5'h4 == index_addr) begin // @[DCache.scala 131:52]
        d2_4 <= 1'h0; // @[DCache.scala 131:52]
      end
    end else if (way2write) begin // @[DCache.scala 132:25]
      d2_4 <= _GEN_1186 | d2_4;
    end
    if (reset) begin // @[DCache.scala 58:26]
      d2_5 <= 1'h0; // @[DCache.scala 58:26]
    end else if (state == 3'h6) begin // @[DCache.scala 130:35]
      if (5'h5 == fence_cnt) begin // @[DCache.scala 130:50]
        d2_5 <= 1'h0; // @[DCache.scala 130:50]
      end
    end else if (update & updateway2) begin // @[DCache.scala 131:36]
      if (5'h5 == index_addr) begin // @[DCache.scala 131:52]
        d2_5 <= 1'h0; // @[DCache.scala 131:52]
      end
    end else if (way2write) begin // @[DCache.scala 132:25]
      d2_5 <= _GEN_1187 | d2_5;
    end
    if (reset) begin // @[DCache.scala 58:26]
      d2_6 <= 1'h0; // @[DCache.scala 58:26]
    end else if (state == 3'h6) begin // @[DCache.scala 130:35]
      if (5'h6 == fence_cnt) begin // @[DCache.scala 130:50]
        d2_6 <= 1'h0; // @[DCache.scala 130:50]
      end
    end else if (update & updateway2) begin // @[DCache.scala 131:36]
      if (5'h6 == index_addr) begin // @[DCache.scala 131:52]
        d2_6 <= 1'h0; // @[DCache.scala 131:52]
      end
    end else if (way2write) begin // @[DCache.scala 132:25]
      d2_6 <= _GEN_1188 | d2_6;
    end
    if (reset) begin // @[DCache.scala 58:26]
      d2_7 <= 1'h0; // @[DCache.scala 58:26]
    end else if (state == 3'h6) begin // @[DCache.scala 130:35]
      if (5'h7 == fence_cnt) begin // @[DCache.scala 130:50]
        d2_7 <= 1'h0; // @[DCache.scala 130:50]
      end
    end else if (update & updateway2) begin // @[DCache.scala 131:36]
      if (5'h7 == index_addr) begin // @[DCache.scala 131:52]
        d2_7 <= 1'h0; // @[DCache.scala 131:52]
      end
    end else if (way2write) begin // @[DCache.scala 132:25]
      d2_7 <= _GEN_1189 | d2_7;
    end
    if (reset) begin // @[DCache.scala 58:26]
      d2_8 <= 1'h0; // @[DCache.scala 58:26]
    end else if (state == 3'h6) begin // @[DCache.scala 130:35]
      if (5'h8 == fence_cnt) begin // @[DCache.scala 130:50]
        d2_8 <= 1'h0; // @[DCache.scala 130:50]
      end
    end else if (update & updateway2) begin // @[DCache.scala 131:36]
      if (5'h8 == index_addr) begin // @[DCache.scala 131:52]
        d2_8 <= 1'h0; // @[DCache.scala 131:52]
      end
    end else if (way2write) begin // @[DCache.scala 132:25]
      d2_8 <= _GEN_1190 | d2_8;
    end
    if (reset) begin // @[DCache.scala 58:26]
      d2_9 <= 1'h0; // @[DCache.scala 58:26]
    end else if (state == 3'h6) begin // @[DCache.scala 130:35]
      if (5'h9 == fence_cnt) begin // @[DCache.scala 130:50]
        d2_9 <= 1'h0; // @[DCache.scala 130:50]
      end
    end else if (update & updateway2) begin // @[DCache.scala 131:36]
      if (5'h9 == index_addr) begin // @[DCache.scala 131:52]
        d2_9 <= 1'h0; // @[DCache.scala 131:52]
      end
    end else if (way2write) begin // @[DCache.scala 132:25]
      d2_9 <= _GEN_1191 | d2_9;
    end
    if (reset) begin // @[DCache.scala 58:26]
      d2_10 <= 1'h0; // @[DCache.scala 58:26]
    end else if (state == 3'h6) begin // @[DCache.scala 130:35]
      if (5'ha == fence_cnt) begin // @[DCache.scala 130:50]
        d2_10 <= 1'h0; // @[DCache.scala 130:50]
      end
    end else if (update & updateway2) begin // @[DCache.scala 131:36]
      if (5'ha == index_addr) begin // @[DCache.scala 131:52]
        d2_10 <= 1'h0; // @[DCache.scala 131:52]
      end
    end else if (way2write) begin // @[DCache.scala 132:25]
      d2_10 <= _GEN_1192 | d2_10;
    end
    if (reset) begin // @[DCache.scala 58:26]
      d2_11 <= 1'h0; // @[DCache.scala 58:26]
    end else if (state == 3'h6) begin // @[DCache.scala 130:35]
      if (5'hb == fence_cnt) begin // @[DCache.scala 130:50]
        d2_11 <= 1'h0; // @[DCache.scala 130:50]
      end
    end else if (update & updateway2) begin // @[DCache.scala 131:36]
      if (5'hb == index_addr) begin // @[DCache.scala 131:52]
        d2_11 <= 1'h0; // @[DCache.scala 131:52]
      end
    end else if (way2write) begin // @[DCache.scala 132:25]
      d2_11 <= _GEN_1193 | d2_11;
    end
    if (reset) begin // @[DCache.scala 58:26]
      d2_12 <= 1'h0; // @[DCache.scala 58:26]
    end else if (state == 3'h6) begin // @[DCache.scala 130:35]
      if (5'hc == fence_cnt) begin // @[DCache.scala 130:50]
        d2_12 <= 1'h0; // @[DCache.scala 130:50]
      end
    end else if (update & updateway2) begin // @[DCache.scala 131:36]
      if (5'hc == index_addr) begin // @[DCache.scala 131:52]
        d2_12 <= 1'h0; // @[DCache.scala 131:52]
      end
    end else if (way2write) begin // @[DCache.scala 132:25]
      d2_12 <= _GEN_1194 | d2_12;
    end
    if (reset) begin // @[DCache.scala 58:26]
      d2_13 <= 1'h0; // @[DCache.scala 58:26]
    end else if (state == 3'h6) begin // @[DCache.scala 130:35]
      if (5'hd == fence_cnt) begin // @[DCache.scala 130:50]
        d2_13 <= 1'h0; // @[DCache.scala 130:50]
      end
    end else if (update & updateway2) begin // @[DCache.scala 131:36]
      if (5'hd == index_addr) begin // @[DCache.scala 131:52]
        d2_13 <= 1'h0; // @[DCache.scala 131:52]
      end
    end else if (way2write) begin // @[DCache.scala 132:25]
      d2_13 <= _GEN_1195 | d2_13;
    end
    if (reset) begin // @[DCache.scala 58:26]
      d2_14 <= 1'h0; // @[DCache.scala 58:26]
    end else if (state == 3'h6) begin // @[DCache.scala 130:35]
      if (5'he == fence_cnt) begin // @[DCache.scala 130:50]
        d2_14 <= 1'h0; // @[DCache.scala 130:50]
      end
    end else if (update & updateway2) begin // @[DCache.scala 131:36]
      if (5'he == index_addr) begin // @[DCache.scala 131:52]
        d2_14 <= 1'h0; // @[DCache.scala 131:52]
      end
    end else if (way2write) begin // @[DCache.scala 132:25]
      d2_14 <= _GEN_1196 | d2_14;
    end
    if (reset) begin // @[DCache.scala 58:26]
      d2_15 <= 1'h0; // @[DCache.scala 58:26]
    end else if (state == 3'h6) begin // @[DCache.scala 130:35]
      if (5'hf == fence_cnt) begin // @[DCache.scala 130:50]
        d2_15 <= 1'h0; // @[DCache.scala 130:50]
      end
    end else if (update & updateway2) begin // @[DCache.scala 131:36]
      if (5'hf == index_addr) begin // @[DCache.scala 131:52]
        d2_15 <= 1'h0; // @[DCache.scala 131:52]
      end
    end else if (way2write) begin // @[DCache.scala 132:25]
      d2_15 <= _GEN_1197 | d2_15;
    end
    if (reset) begin // @[DCache.scala 58:26]
      d2_16 <= 1'h0; // @[DCache.scala 58:26]
    end else if (state == 3'h6) begin // @[DCache.scala 130:35]
      if (5'h10 == fence_cnt) begin // @[DCache.scala 130:50]
        d2_16 <= 1'h0; // @[DCache.scala 130:50]
      end
    end else if (update & updateway2) begin // @[DCache.scala 131:36]
      if (5'h10 == index_addr) begin // @[DCache.scala 131:52]
        d2_16 <= 1'h0; // @[DCache.scala 131:52]
      end
    end else if (way2write) begin // @[DCache.scala 132:25]
      d2_16 <= _GEN_1198 | d2_16;
    end
    if (reset) begin // @[DCache.scala 58:26]
      d2_17 <= 1'h0; // @[DCache.scala 58:26]
    end else if (state == 3'h6) begin // @[DCache.scala 130:35]
      if (5'h11 == fence_cnt) begin // @[DCache.scala 130:50]
        d2_17 <= 1'h0; // @[DCache.scala 130:50]
      end
    end else if (update & updateway2) begin // @[DCache.scala 131:36]
      if (5'h11 == index_addr) begin // @[DCache.scala 131:52]
        d2_17 <= 1'h0; // @[DCache.scala 131:52]
      end
    end else if (way2write) begin // @[DCache.scala 132:25]
      d2_17 <= _GEN_1199 | d2_17;
    end
    if (reset) begin // @[DCache.scala 58:26]
      d2_18 <= 1'h0; // @[DCache.scala 58:26]
    end else if (state == 3'h6) begin // @[DCache.scala 130:35]
      if (5'h12 == fence_cnt) begin // @[DCache.scala 130:50]
        d2_18 <= 1'h0; // @[DCache.scala 130:50]
      end
    end else if (update & updateway2) begin // @[DCache.scala 131:36]
      if (5'h12 == index_addr) begin // @[DCache.scala 131:52]
        d2_18 <= 1'h0; // @[DCache.scala 131:52]
      end
    end else if (way2write) begin // @[DCache.scala 132:25]
      d2_18 <= _GEN_1200 | d2_18;
    end
    if (reset) begin // @[DCache.scala 58:26]
      d2_19 <= 1'h0; // @[DCache.scala 58:26]
    end else if (state == 3'h6) begin // @[DCache.scala 130:35]
      if (5'h13 == fence_cnt) begin // @[DCache.scala 130:50]
        d2_19 <= 1'h0; // @[DCache.scala 130:50]
      end
    end else if (update & updateway2) begin // @[DCache.scala 131:36]
      if (5'h13 == index_addr) begin // @[DCache.scala 131:52]
        d2_19 <= 1'h0; // @[DCache.scala 131:52]
      end
    end else if (way2write) begin // @[DCache.scala 132:25]
      d2_19 <= _GEN_1201 | d2_19;
    end
    if (reset) begin // @[DCache.scala 58:26]
      d2_20 <= 1'h0; // @[DCache.scala 58:26]
    end else if (state == 3'h6) begin // @[DCache.scala 130:35]
      if (5'h14 == fence_cnt) begin // @[DCache.scala 130:50]
        d2_20 <= 1'h0; // @[DCache.scala 130:50]
      end
    end else if (update & updateway2) begin // @[DCache.scala 131:36]
      if (5'h14 == index_addr) begin // @[DCache.scala 131:52]
        d2_20 <= 1'h0; // @[DCache.scala 131:52]
      end
    end else if (way2write) begin // @[DCache.scala 132:25]
      d2_20 <= _GEN_1202 | d2_20;
    end
    if (reset) begin // @[DCache.scala 58:26]
      d2_21 <= 1'h0; // @[DCache.scala 58:26]
    end else if (state == 3'h6) begin // @[DCache.scala 130:35]
      if (5'h15 == fence_cnt) begin // @[DCache.scala 130:50]
        d2_21 <= 1'h0; // @[DCache.scala 130:50]
      end
    end else if (update & updateway2) begin // @[DCache.scala 131:36]
      if (5'h15 == index_addr) begin // @[DCache.scala 131:52]
        d2_21 <= 1'h0; // @[DCache.scala 131:52]
      end
    end else if (way2write) begin // @[DCache.scala 132:25]
      d2_21 <= _GEN_1203 | d2_21;
    end
    if (reset) begin // @[DCache.scala 58:26]
      d2_22 <= 1'h0; // @[DCache.scala 58:26]
    end else if (state == 3'h6) begin // @[DCache.scala 130:35]
      if (5'h16 == fence_cnt) begin // @[DCache.scala 130:50]
        d2_22 <= 1'h0; // @[DCache.scala 130:50]
      end
    end else if (update & updateway2) begin // @[DCache.scala 131:36]
      if (5'h16 == index_addr) begin // @[DCache.scala 131:52]
        d2_22 <= 1'h0; // @[DCache.scala 131:52]
      end
    end else if (way2write) begin // @[DCache.scala 132:25]
      d2_22 <= _GEN_1204 | d2_22;
    end
    if (reset) begin // @[DCache.scala 58:26]
      d2_23 <= 1'h0; // @[DCache.scala 58:26]
    end else if (state == 3'h6) begin // @[DCache.scala 130:35]
      if (5'h17 == fence_cnt) begin // @[DCache.scala 130:50]
        d2_23 <= 1'h0; // @[DCache.scala 130:50]
      end
    end else if (update & updateway2) begin // @[DCache.scala 131:36]
      if (5'h17 == index_addr) begin // @[DCache.scala 131:52]
        d2_23 <= 1'h0; // @[DCache.scala 131:52]
      end
    end else if (way2write) begin // @[DCache.scala 132:25]
      d2_23 <= _GEN_1205 | d2_23;
    end
    if (reset) begin // @[DCache.scala 58:26]
      d2_24 <= 1'h0; // @[DCache.scala 58:26]
    end else if (state == 3'h6) begin // @[DCache.scala 130:35]
      if (5'h18 == fence_cnt) begin // @[DCache.scala 130:50]
        d2_24 <= 1'h0; // @[DCache.scala 130:50]
      end
    end else if (update & updateway2) begin // @[DCache.scala 131:36]
      if (5'h18 == index_addr) begin // @[DCache.scala 131:52]
        d2_24 <= 1'h0; // @[DCache.scala 131:52]
      end
    end else if (way2write) begin // @[DCache.scala 132:25]
      d2_24 <= _GEN_1206 | d2_24;
    end
    if (reset) begin // @[DCache.scala 58:26]
      d2_25 <= 1'h0; // @[DCache.scala 58:26]
    end else if (state == 3'h6) begin // @[DCache.scala 130:35]
      if (5'h19 == fence_cnt) begin // @[DCache.scala 130:50]
        d2_25 <= 1'h0; // @[DCache.scala 130:50]
      end
    end else if (update & updateway2) begin // @[DCache.scala 131:36]
      if (5'h19 == index_addr) begin // @[DCache.scala 131:52]
        d2_25 <= 1'h0; // @[DCache.scala 131:52]
      end
    end else if (way2write) begin // @[DCache.scala 132:25]
      d2_25 <= _GEN_1207 | d2_25;
    end
    if (reset) begin // @[DCache.scala 58:26]
      d2_26 <= 1'h0; // @[DCache.scala 58:26]
    end else if (state == 3'h6) begin // @[DCache.scala 130:35]
      if (5'h1a == fence_cnt) begin // @[DCache.scala 130:50]
        d2_26 <= 1'h0; // @[DCache.scala 130:50]
      end
    end else if (update & updateway2) begin // @[DCache.scala 131:36]
      if (5'h1a == index_addr) begin // @[DCache.scala 131:52]
        d2_26 <= 1'h0; // @[DCache.scala 131:52]
      end
    end else if (way2write) begin // @[DCache.scala 132:25]
      d2_26 <= _GEN_1208 | d2_26;
    end
    if (reset) begin // @[DCache.scala 58:26]
      d2_27 <= 1'h0; // @[DCache.scala 58:26]
    end else if (state == 3'h6) begin // @[DCache.scala 130:35]
      if (5'h1b == fence_cnt) begin // @[DCache.scala 130:50]
        d2_27 <= 1'h0; // @[DCache.scala 130:50]
      end
    end else if (update & updateway2) begin // @[DCache.scala 131:36]
      if (5'h1b == index_addr) begin // @[DCache.scala 131:52]
        d2_27 <= 1'h0; // @[DCache.scala 131:52]
      end
    end else if (way2write) begin // @[DCache.scala 132:25]
      d2_27 <= _GEN_1209 | d2_27;
    end
    if (reset) begin // @[DCache.scala 58:26]
      d2_28 <= 1'h0; // @[DCache.scala 58:26]
    end else if (state == 3'h6) begin // @[DCache.scala 130:35]
      if (5'h1c == fence_cnt) begin // @[DCache.scala 130:50]
        d2_28 <= 1'h0; // @[DCache.scala 130:50]
      end
    end else if (update & updateway2) begin // @[DCache.scala 131:36]
      if (5'h1c == index_addr) begin // @[DCache.scala 131:52]
        d2_28 <= 1'h0; // @[DCache.scala 131:52]
      end
    end else if (way2write) begin // @[DCache.scala 132:25]
      d2_28 <= _GEN_1210 | d2_28;
    end
    if (reset) begin // @[DCache.scala 58:26]
      d2_29 <= 1'h0; // @[DCache.scala 58:26]
    end else if (state == 3'h6) begin // @[DCache.scala 130:35]
      if (5'h1d == fence_cnt) begin // @[DCache.scala 130:50]
        d2_29 <= 1'h0; // @[DCache.scala 130:50]
      end
    end else if (update & updateway2) begin // @[DCache.scala 131:36]
      if (5'h1d == index_addr) begin // @[DCache.scala 131:52]
        d2_29 <= 1'h0; // @[DCache.scala 131:52]
      end
    end else if (way2write) begin // @[DCache.scala 132:25]
      d2_29 <= _GEN_1211 | d2_29;
    end
    if (reset) begin // @[DCache.scala 58:26]
      d2_30 <= 1'h0; // @[DCache.scala 58:26]
    end else if (state == 3'h6) begin // @[DCache.scala 130:35]
      if (5'h1e == fence_cnt) begin // @[DCache.scala 130:50]
        d2_30 <= 1'h0; // @[DCache.scala 130:50]
      end
    end else if (update & updateway2) begin // @[DCache.scala 131:36]
      if (5'h1e == index_addr) begin // @[DCache.scala 131:52]
        d2_30 <= 1'h0; // @[DCache.scala 131:52]
      end
    end else if (way2write) begin // @[DCache.scala 132:25]
      d2_30 <= _GEN_1212 | d2_30;
    end
    if (reset) begin // @[DCache.scala 58:26]
      d2_31 <= 1'h0; // @[DCache.scala 58:26]
    end else if (state == 3'h6) begin // @[DCache.scala 130:35]
      if (5'h1f == fence_cnt) begin // @[DCache.scala 130:50]
        d2_31 <= 1'h0; // @[DCache.scala 130:50]
      end
    end else if (update & updateway2) begin // @[DCache.scala 131:36]
      if (5'h1f == index_addr) begin // @[DCache.scala 131:52]
        d2_31 <= 1'h0; // @[DCache.scala 131:52]
      end
    end else if (way2write) begin // @[DCache.scala 132:25]
      d2_31 <= _GEN_1213 | d2_31;
    end
    if (reset) begin // @[DCache.scala 59:26]
      age2_0 <= 1'h0; // @[DCache.scala 59:26]
    end else if (5'h0 == index_addr) begin // @[DCache.scala 82:22]
      if (_age1_T) begin // @[DCache.scala 82:28]
        age2_0 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 82:28]
        age2_0 <= age2_31; // @[DCache.scala 82:28]
      end else begin
        age2_0 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 59:26]
      age2_1 <= 1'h0; // @[DCache.scala 59:26]
    end else if (5'h1 == index_addr) begin // @[DCache.scala 82:22]
      if (_age1_T) begin // @[DCache.scala 82:28]
        age2_1 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 82:28]
        age2_1 <= age2_31; // @[DCache.scala 82:28]
      end else begin
        age2_1 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 59:26]
      age2_2 <= 1'h0; // @[DCache.scala 59:26]
    end else if (5'h2 == index_addr) begin // @[DCache.scala 82:22]
      if (_age1_T) begin // @[DCache.scala 82:28]
        age2_2 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 82:28]
        age2_2 <= age2_31; // @[DCache.scala 82:28]
      end else begin
        age2_2 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 59:26]
      age2_3 <= 1'h0; // @[DCache.scala 59:26]
    end else if (5'h3 == index_addr) begin // @[DCache.scala 82:22]
      if (_age1_T) begin // @[DCache.scala 82:28]
        age2_3 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 82:28]
        age2_3 <= age2_31; // @[DCache.scala 82:28]
      end else begin
        age2_3 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 59:26]
      age2_4 <= 1'h0; // @[DCache.scala 59:26]
    end else if (5'h4 == index_addr) begin // @[DCache.scala 82:22]
      if (_age1_T) begin // @[DCache.scala 82:28]
        age2_4 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 82:28]
        age2_4 <= age2_31; // @[DCache.scala 82:28]
      end else begin
        age2_4 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 59:26]
      age2_5 <= 1'h0; // @[DCache.scala 59:26]
    end else if (5'h5 == index_addr) begin // @[DCache.scala 82:22]
      if (_age1_T) begin // @[DCache.scala 82:28]
        age2_5 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 82:28]
        age2_5 <= age2_31; // @[DCache.scala 82:28]
      end else begin
        age2_5 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 59:26]
      age2_6 <= 1'h0; // @[DCache.scala 59:26]
    end else if (5'h6 == index_addr) begin // @[DCache.scala 82:22]
      if (_age1_T) begin // @[DCache.scala 82:28]
        age2_6 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 82:28]
        age2_6 <= age2_31; // @[DCache.scala 82:28]
      end else begin
        age2_6 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 59:26]
      age2_7 <= 1'h0; // @[DCache.scala 59:26]
    end else if (5'h7 == index_addr) begin // @[DCache.scala 82:22]
      if (_age1_T) begin // @[DCache.scala 82:28]
        age2_7 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 82:28]
        age2_7 <= age2_31; // @[DCache.scala 82:28]
      end else begin
        age2_7 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 59:26]
      age2_8 <= 1'h0; // @[DCache.scala 59:26]
    end else if (5'h8 == index_addr) begin // @[DCache.scala 82:22]
      if (_age1_T) begin // @[DCache.scala 82:28]
        age2_8 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 82:28]
        age2_8 <= age2_31; // @[DCache.scala 82:28]
      end else begin
        age2_8 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 59:26]
      age2_9 <= 1'h0; // @[DCache.scala 59:26]
    end else if (5'h9 == index_addr) begin // @[DCache.scala 82:22]
      if (_age1_T) begin // @[DCache.scala 82:28]
        age2_9 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 82:28]
        age2_9 <= age2_31; // @[DCache.scala 82:28]
      end else begin
        age2_9 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 59:26]
      age2_10 <= 1'h0; // @[DCache.scala 59:26]
    end else if (5'ha == index_addr) begin // @[DCache.scala 82:22]
      if (_age1_T) begin // @[DCache.scala 82:28]
        age2_10 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 82:28]
        age2_10 <= age2_31; // @[DCache.scala 82:28]
      end else begin
        age2_10 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 59:26]
      age2_11 <= 1'h0; // @[DCache.scala 59:26]
    end else if (5'hb == index_addr) begin // @[DCache.scala 82:22]
      if (_age1_T) begin // @[DCache.scala 82:28]
        age2_11 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 82:28]
        age2_11 <= age2_31; // @[DCache.scala 82:28]
      end else begin
        age2_11 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 59:26]
      age2_12 <= 1'h0; // @[DCache.scala 59:26]
    end else if (5'hc == index_addr) begin // @[DCache.scala 82:22]
      if (_age1_T) begin // @[DCache.scala 82:28]
        age2_12 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 82:28]
        age2_12 <= age2_31; // @[DCache.scala 82:28]
      end else begin
        age2_12 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 59:26]
      age2_13 <= 1'h0; // @[DCache.scala 59:26]
    end else if (5'hd == index_addr) begin // @[DCache.scala 82:22]
      if (_age1_T) begin // @[DCache.scala 82:28]
        age2_13 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 82:28]
        age2_13 <= age2_31; // @[DCache.scala 82:28]
      end else begin
        age2_13 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 59:26]
      age2_14 <= 1'h0; // @[DCache.scala 59:26]
    end else if (5'he == index_addr) begin // @[DCache.scala 82:22]
      if (_age1_T) begin // @[DCache.scala 82:28]
        age2_14 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 82:28]
        age2_14 <= age2_31; // @[DCache.scala 82:28]
      end else begin
        age2_14 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 59:26]
      age2_15 <= 1'h0; // @[DCache.scala 59:26]
    end else if (5'hf == index_addr) begin // @[DCache.scala 82:22]
      if (_age1_T) begin // @[DCache.scala 82:28]
        age2_15 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 82:28]
        age2_15 <= age2_31; // @[DCache.scala 82:28]
      end else begin
        age2_15 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 59:26]
      age2_16 <= 1'h0; // @[DCache.scala 59:26]
    end else if (5'h10 == index_addr) begin // @[DCache.scala 82:22]
      if (_age1_T) begin // @[DCache.scala 82:28]
        age2_16 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 82:28]
        age2_16 <= age2_31; // @[DCache.scala 82:28]
      end else begin
        age2_16 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 59:26]
      age2_17 <= 1'h0; // @[DCache.scala 59:26]
    end else if (5'h11 == index_addr) begin // @[DCache.scala 82:22]
      if (_age1_T) begin // @[DCache.scala 82:28]
        age2_17 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 82:28]
        age2_17 <= age2_31; // @[DCache.scala 82:28]
      end else begin
        age2_17 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 59:26]
      age2_18 <= 1'h0; // @[DCache.scala 59:26]
    end else if (5'h12 == index_addr) begin // @[DCache.scala 82:22]
      if (_age1_T) begin // @[DCache.scala 82:28]
        age2_18 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 82:28]
        age2_18 <= age2_31; // @[DCache.scala 82:28]
      end else begin
        age2_18 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 59:26]
      age2_19 <= 1'h0; // @[DCache.scala 59:26]
    end else if (5'h13 == index_addr) begin // @[DCache.scala 82:22]
      if (_age1_T) begin // @[DCache.scala 82:28]
        age2_19 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 82:28]
        age2_19 <= age2_31; // @[DCache.scala 82:28]
      end else begin
        age2_19 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 59:26]
      age2_20 <= 1'h0; // @[DCache.scala 59:26]
    end else if (5'h14 == index_addr) begin // @[DCache.scala 82:22]
      if (_age1_T) begin // @[DCache.scala 82:28]
        age2_20 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 82:28]
        age2_20 <= age2_31; // @[DCache.scala 82:28]
      end else begin
        age2_20 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 59:26]
      age2_21 <= 1'h0; // @[DCache.scala 59:26]
    end else if (5'h15 == index_addr) begin // @[DCache.scala 82:22]
      if (_age1_T) begin // @[DCache.scala 82:28]
        age2_21 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 82:28]
        age2_21 <= age2_31; // @[DCache.scala 82:28]
      end else begin
        age2_21 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 59:26]
      age2_22 <= 1'h0; // @[DCache.scala 59:26]
    end else if (5'h16 == index_addr) begin // @[DCache.scala 82:22]
      if (_age1_T) begin // @[DCache.scala 82:28]
        age2_22 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 82:28]
        age2_22 <= age2_31; // @[DCache.scala 82:28]
      end else begin
        age2_22 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 59:26]
      age2_23 <= 1'h0; // @[DCache.scala 59:26]
    end else if (5'h17 == index_addr) begin // @[DCache.scala 82:22]
      if (_age1_T) begin // @[DCache.scala 82:28]
        age2_23 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 82:28]
        age2_23 <= age2_31; // @[DCache.scala 82:28]
      end else begin
        age2_23 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 59:26]
      age2_24 <= 1'h0; // @[DCache.scala 59:26]
    end else if (5'h18 == index_addr) begin // @[DCache.scala 82:22]
      if (_age1_T) begin // @[DCache.scala 82:28]
        age2_24 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 82:28]
        age2_24 <= age2_31; // @[DCache.scala 82:28]
      end else begin
        age2_24 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 59:26]
      age2_25 <= 1'h0; // @[DCache.scala 59:26]
    end else if (5'h19 == index_addr) begin // @[DCache.scala 82:22]
      if (_age1_T) begin // @[DCache.scala 82:28]
        age2_25 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 82:28]
        age2_25 <= age2_31; // @[DCache.scala 82:28]
      end else begin
        age2_25 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 59:26]
      age2_26 <= 1'h0; // @[DCache.scala 59:26]
    end else if (5'h1a == index_addr) begin // @[DCache.scala 82:22]
      if (_age1_T) begin // @[DCache.scala 82:28]
        age2_26 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 82:28]
        age2_26 <= age2_31; // @[DCache.scala 82:28]
      end else begin
        age2_26 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 59:26]
      age2_27 <= 1'h0; // @[DCache.scala 59:26]
    end else if (5'h1b == index_addr) begin // @[DCache.scala 82:22]
      if (_age1_T) begin // @[DCache.scala 82:28]
        age2_27 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 82:28]
        age2_27 <= age2_31; // @[DCache.scala 82:28]
      end else begin
        age2_27 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 59:26]
      age2_28 <= 1'h0; // @[DCache.scala 59:26]
    end else if (5'h1c == index_addr) begin // @[DCache.scala 82:22]
      if (_age1_T) begin // @[DCache.scala 82:28]
        age2_28 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 82:28]
        age2_28 <= age2_31; // @[DCache.scala 82:28]
      end else begin
        age2_28 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 59:26]
      age2_29 <= 1'h0; // @[DCache.scala 59:26]
    end else if (5'h1d == index_addr) begin // @[DCache.scala 82:22]
      if (_age1_T) begin // @[DCache.scala 82:28]
        age2_29 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 82:28]
        age2_29 <= age2_31; // @[DCache.scala 82:28]
      end else begin
        age2_29 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 59:26]
      age2_30 <= 1'h0; // @[DCache.scala 59:26]
    end else if (5'h1e == index_addr) begin // @[DCache.scala 82:22]
      if (_age1_T) begin // @[DCache.scala 82:28]
        age2_30 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 82:28]
        age2_30 <= age2_31; // @[DCache.scala 82:28]
      end else begin
        age2_30 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 59:26]
      age2_31 <= 1'h0; // @[DCache.scala 59:26]
    end else if (5'h1f == index_addr) begin // @[DCache.scala 82:22]
      if (_age1_T) begin // @[DCache.scala 82:28]
        age2_31 <= hit2;
      end else if (!(5'h1f == index_addr)) begin // @[DCache.scala 82:28]
        age2_31 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 60:26]
      tag2_0 <= 53'h0; // @[DCache.scala 60:26]
    end else if (5'h0 == index_addr) begin // @[DCache.scala 147:26]
      if (_T_22) begin // @[DCache.scala 147:32]
        tag2_0 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 64:28]
        tag2_0 <= tag2_31; // @[DCache.scala 64:28]
      end else begin
        tag2_0 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 60:26]
      tag2_1 <= 53'h0; // @[DCache.scala 60:26]
    end else if (5'h1 == index_addr) begin // @[DCache.scala 147:26]
      if (_T_22) begin // @[DCache.scala 147:32]
        tag2_1 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 64:28]
        tag2_1 <= tag2_31; // @[DCache.scala 64:28]
      end else begin
        tag2_1 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 60:26]
      tag2_2 <= 53'h0; // @[DCache.scala 60:26]
    end else if (5'h2 == index_addr) begin // @[DCache.scala 147:26]
      if (_T_22) begin // @[DCache.scala 147:32]
        tag2_2 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 64:28]
        tag2_2 <= tag2_31; // @[DCache.scala 64:28]
      end else begin
        tag2_2 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 60:26]
      tag2_3 <= 53'h0; // @[DCache.scala 60:26]
    end else if (5'h3 == index_addr) begin // @[DCache.scala 147:26]
      if (_T_22) begin // @[DCache.scala 147:32]
        tag2_3 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 64:28]
        tag2_3 <= tag2_31; // @[DCache.scala 64:28]
      end else begin
        tag2_3 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 60:26]
      tag2_4 <= 53'h0; // @[DCache.scala 60:26]
    end else if (5'h4 == index_addr) begin // @[DCache.scala 147:26]
      if (_T_22) begin // @[DCache.scala 147:32]
        tag2_4 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 64:28]
        tag2_4 <= tag2_31; // @[DCache.scala 64:28]
      end else begin
        tag2_4 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 60:26]
      tag2_5 <= 53'h0; // @[DCache.scala 60:26]
    end else if (5'h5 == index_addr) begin // @[DCache.scala 147:26]
      if (_T_22) begin // @[DCache.scala 147:32]
        tag2_5 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 64:28]
        tag2_5 <= tag2_31; // @[DCache.scala 64:28]
      end else begin
        tag2_5 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 60:26]
      tag2_6 <= 53'h0; // @[DCache.scala 60:26]
    end else if (5'h6 == index_addr) begin // @[DCache.scala 147:26]
      if (_T_22) begin // @[DCache.scala 147:32]
        tag2_6 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 64:28]
        tag2_6 <= tag2_31; // @[DCache.scala 64:28]
      end else begin
        tag2_6 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 60:26]
      tag2_7 <= 53'h0; // @[DCache.scala 60:26]
    end else if (5'h7 == index_addr) begin // @[DCache.scala 147:26]
      if (_T_22) begin // @[DCache.scala 147:32]
        tag2_7 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 64:28]
        tag2_7 <= tag2_31; // @[DCache.scala 64:28]
      end else begin
        tag2_7 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 60:26]
      tag2_8 <= 53'h0; // @[DCache.scala 60:26]
    end else if (5'h8 == index_addr) begin // @[DCache.scala 147:26]
      if (_T_22) begin // @[DCache.scala 147:32]
        tag2_8 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 64:28]
        tag2_8 <= tag2_31; // @[DCache.scala 64:28]
      end else begin
        tag2_8 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 60:26]
      tag2_9 <= 53'h0; // @[DCache.scala 60:26]
    end else if (5'h9 == index_addr) begin // @[DCache.scala 147:26]
      if (_T_22) begin // @[DCache.scala 147:32]
        tag2_9 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 64:28]
        tag2_9 <= tag2_31; // @[DCache.scala 64:28]
      end else begin
        tag2_9 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 60:26]
      tag2_10 <= 53'h0; // @[DCache.scala 60:26]
    end else if (5'ha == index_addr) begin // @[DCache.scala 147:26]
      if (_T_22) begin // @[DCache.scala 147:32]
        tag2_10 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 64:28]
        tag2_10 <= tag2_31; // @[DCache.scala 64:28]
      end else begin
        tag2_10 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 60:26]
      tag2_11 <= 53'h0; // @[DCache.scala 60:26]
    end else if (5'hb == index_addr) begin // @[DCache.scala 147:26]
      if (_T_22) begin // @[DCache.scala 147:32]
        tag2_11 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 64:28]
        tag2_11 <= tag2_31; // @[DCache.scala 64:28]
      end else begin
        tag2_11 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 60:26]
      tag2_12 <= 53'h0; // @[DCache.scala 60:26]
    end else if (5'hc == index_addr) begin // @[DCache.scala 147:26]
      if (_T_22) begin // @[DCache.scala 147:32]
        tag2_12 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 64:28]
        tag2_12 <= tag2_31; // @[DCache.scala 64:28]
      end else begin
        tag2_12 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 60:26]
      tag2_13 <= 53'h0; // @[DCache.scala 60:26]
    end else if (5'hd == index_addr) begin // @[DCache.scala 147:26]
      if (_T_22) begin // @[DCache.scala 147:32]
        tag2_13 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 64:28]
        tag2_13 <= tag2_31; // @[DCache.scala 64:28]
      end else begin
        tag2_13 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 60:26]
      tag2_14 <= 53'h0; // @[DCache.scala 60:26]
    end else if (5'he == index_addr) begin // @[DCache.scala 147:26]
      if (_T_22) begin // @[DCache.scala 147:32]
        tag2_14 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 64:28]
        tag2_14 <= tag2_31; // @[DCache.scala 64:28]
      end else begin
        tag2_14 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 60:26]
      tag2_15 <= 53'h0; // @[DCache.scala 60:26]
    end else if (5'hf == index_addr) begin // @[DCache.scala 147:26]
      if (_T_22) begin // @[DCache.scala 147:32]
        tag2_15 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 64:28]
        tag2_15 <= tag2_31; // @[DCache.scala 64:28]
      end else begin
        tag2_15 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 60:26]
      tag2_16 <= 53'h0; // @[DCache.scala 60:26]
    end else if (5'h10 == index_addr) begin // @[DCache.scala 147:26]
      if (_T_22) begin // @[DCache.scala 147:32]
        tag2_16 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 64:28]
        tag2_16 <= tag2_31; // @[DCache.scala 64:28]
      end else begin
        tag2_16 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 60:26]
      tag2_17 <= 53'h0; // @[DCache.scala 60:26]
    end else if (5'h11 == index_addr) begin // @[DCache.scala 147:26]
      if (_T_22) begin // @[DCache.scala 147:32]
        tag2_17 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 64:28]
        tag2_17 <= tag2_31; // @[DCache.scala 64:28]
      end else begin
        tag2_17 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 60:26]
      tag2_18 <= 53'h0; // @[DCache.scala 60:26]
    end else if (5'h12 == index_addr) begin // @[DCache.scala 147:26]
      if (_T_22) begin // @[DCache.scala 147:32]
        tag2_18 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 64:28]
        tag2_18 <= tag2_31; // @[DCache.scala 64:28]
      end else begin
        tag2_18 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 60:26]
      tag2_19 <= 53'h0; // @[DCache.scala 60:26]
    end else if (5'h13 == index_addr) begin // @[DCache.scala 147:26]
      if (_T_22) begin // @[DCache.scala 147:32]
        tag2_19 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 64:28]
        tag2_19 <= tag2_31; // @[DCache.scala 64:28]
      end else begin
        tag2_19 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 60:26]
      tag2_20 <= 53'h0; // @[DCache.scala 60:26]
    end else if (5'h14 == index_addr) begin // @[DCache.scala 147:26]
      if (_T_22) begin // @[DCache.scala 147:32]
        tag2_20 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 64:28]
        tag2_20 <= tag2_31; // @[DCache.scala 64:28]
      end else begin
        tag2_20 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 60:26]
      tag2_21 <= 53'h0; // @[DCache.scala 60:26]
    end else if (5'h15 == index_addr) begin // @[DCache.scala 147:26]
      if (_T_22) begin // @[DCache.scala 147:32]
        tag2_21 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 64:28]
        tag2_21 <= tag2_31; // @[DCache.scala 64:28]
      end else begin
        tag2_21 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 60:26]
      tag2_22 <= 53'h0; // @[DCache.scala 60:26]
    end else if (5'h16 == index_addr) begin // @[DCache.scala 147:26]
      if (_T_22) begin // @[DCache.scala 147:32]
        tag2_22 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 64:28]
        tag2_22 <= tag2_31; // @[DCache.scala 64:28]
      end else begin
        tag2_22 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 60:26]
      tag2_23 <= 53'h0; // @[DCache.scala 60:26]
    end else if (5'h17 == index_addr) begin // @[DCache.scala 147:26]
      if (_T_22) begin // @[DCache.scala 147:32]
        tag2_23 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 64:28]
        tag2_23 <= tag2_31; // @[DCache.scala 64:28]
      end else begin
        tag2_23 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 60:26]
      tag2_24 <= 53'h0; // @[DCache.scala 60:26]
    end else if (5'h18 == index_addr) begin // @[DCache.scala 147:26]
      if (_T_22) begin // @[DCache.scala 147:32]
        tag2_24 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 64:28]
        tag2_24 <= tag2_31; // @[DCache.scala 64:28]
      end else begin
        tag2_24 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 60:26]
      tag2_25 <= 53'h0; // @[DCache.scala 60:26]
    end else if (5'h19 == index_addr) begin // @[DCache.scala 147:26]
      if (_T_22) begin // @[DCache.scala 147:32]
        tag2_25 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 64:28]
        tag2_25 <= tag2_31; // @[DCache.scala 64:28]
      end else begin
        tag2_25 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 60:26]
      tag2_26 <= 53'h0; // @[DCache.scala 60:26]
    end else if (5'h1a == index_addr) begin // @[DCache.scala 147:26]
      if (_T_22) begin // @[DCache.scala 147:32]
        tag2_26 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 64:28]
        tag2_26 <= tag2_31; // @[DCache.scala 64:28]
      end else begin
        tag2_26 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 60:26]
      tag2_27 <= 53'h0; // @[DCache.scala 60:26]
    end else if (5'h1b == index_addr) begin // @[DCache.scala 147:26]
      if (_T_22) begin // @[DCache.scala 147:32]
        tag2_27 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 64:28]
        tag2_27 <= tag2_31; // @[DCache.scala 64:28]
      end else begin
        tag2_27 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 60:26]
      tag2_28 <= 53'h0; // @[DCache.scala 60:26]
    end else if (5'h1c == index_addr) begin // @[DCache.scala 147:26]
      if (_T_22) begin // @[DCache.scala 147:32]
        tag2_28 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 64:28]
        tag2_28 <= tag2_31; // @[DCache.scala 64:28]
      end else begin
        tag2_28 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 60:26]
      tag2_29 <= 53'h0; // @[DCache.scala 60:26]
    end else if (5'h1d == index_addr) begin // @[DCache.scala 147:26]
      if (_T_22) begin // @[DCache.scala 147:32]
        tag2_29 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 64:28]
        tag2_29 <= tag2_31; // @[DCache.scala 64:28]
      end else begin
        tag2_29 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 60:26]
      tag2_30 <= 53'h0; // @[DCache.scala 60:26]
    end else if (5'h1e == index_addr) begin // @[DCache.scala 147:26]
      if (_T_22) begin // @[DCache.scala 147:32]
        tag2_30 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 64:28]
        tag2_30 <= tag2_31; // @[DCache.scala 64:28]
      end else begin
        tag2_30 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 60:26]
      tag2_31 <= 53'h0; // @[DCache.scala 60:26]
    end else if (5'h1f == index_addr) begin // @[DCache.scala 147:26]
      if (_T_22) begin // @[DCache.scala 147:32]
        tag2_31 <= tag_addr;
      end else if (!(5'h1f == index_addr)) begin // @[DCache.scala 64:28]
        tag2_31 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 61:26]
      block2_0 <= 512'h0; // @[DCache.scala 61:26]
    end else if (5'h0 == index_addr) begin // @[DCache.scala 146:26]
      if (_T_22) begin // @[DCache.scala 146:32]
        block2_0 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 146:72]
        block2_0 <= block2_after_write;
      end else begin
        block2_0 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 61:26]
      block2_1 <= 512'h0; // @[DCache.scala 61:26]
    end else if (5'h1 == index_addr) begin // @[DCache.scala 146:26]
      if (_T_22) begin // @[DCache.scala 146:32]
        block2_1 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 146:72]
        block2_1 <= block2_after_write;
      end else begin
        block2_1 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 61:26]
      block2_2 <= 512'h0; // @[DCache.scala 61:26]
    end else if (5'h2 == index_addr) begin // @[DCache.scala 146:26]
      if (_T_22) begin // @[DCache.scala 146:32]
        block2_2 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 146:72]
        block2_2 <= block2_after_write;
      end else begin
        block2_2 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 61:26]
      block2_3 <= 512'h0; // @[DCache.scala 61:26]
    end else if (5'h3 == index_addr) begin // @[DCache.scala 146:26]
      if (_T_22) begin // @[DCache.scala 146:32]
        block2_3 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 146:72]
        block2_3 <= block2_after_write;
      end else begin
        block2_3 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 61:26]
      block2_4 <= 512'h0; // @[DCache.scala 61:26]
    end else if (5'h4 == index_addr) begin // @[DCache.scala 146:26]
      if (_T_22) begin // @[DCache.scala 146:32]
        block2_4 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 146:72]
        block2_4 <= block2_after_write;
      end else begin
        block2_4 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 61:26]
      block2_5 <= 512'h0; // @[DCache.scala 61:26]
    end else if (5'h5 == index_addr) begin // @[DCache.scala 146:26]
      if (_T_22) begin // @[DCache.scala 146:32]
        block2_5 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 146:72]
        block2_5 <= block2_after_write;
      end else begin
        block2_5 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 61:26]
      block2_6 <= 512'h0; // @[DCache.scala 61:26]
    end else if (5'h6 == index_addr) begin // @[DCache.scala 146:26]
      if (_T_22) begin // @[DCache.scala 146:32]
        block2_6 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 146:72]
        block2_6 <= block2_after_write;
      end else begin
        block2_6 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 61:26]
      block2_7 <= 512'h0; // @[DCache.scala 61:26]
    end else if (5'h7 == index_addr) begin // @[DCache.scala 146:26]
      if (_T_22) begin // @[DCache.scala 146:32]
        block2_7 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 146:72]
        block2_7 <= block2_after_write;
      end else begin
        block2_7 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 61:26]
      block2_8 <= 512'h0; // @[DCache.scala 61:26]
    end else if (5'h8 == index_addr) begin // @[DCache.scala 146:26]
      if (_T_22) begin // @[DCache.scala 146:32]
        block2_8 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 146:72]
        block2_8 <= block2_after_write;
      end else begin
        block2_8 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 61:26]
      block2_9 <= 512'h0; // @[DCache.scala 61:26]
    end else if (5'h9 == index_addr) begin // @[DCache.scala 146:26]
      if (_T_22) begin // @[DCache.scala 146:32]
        block2_9 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 146:72]
        block2_9 <= block2_after_write;
      end else begin
        block2_9 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 61:26]
      block2_10 <= 512'h0; // @[DCache.scala 61:26]
    end else if (5'ha == index_addr) begin // @[DCache.scala 146:26]
      if (_T_22) begin // @[DCache.scala 146:32]
        block2_10 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 146:72]
        block2_10 <= block2_after_write;
      end else begin
        block2_10 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 61:26]
      block2_11 <= 512'h0; // @[DCache.scala 61:26]
    end else if (5'hb == index_addr) begin // @[DCache.scala 146:26]
      if (_T_22) begin // @[DCache.scala 146:32]
        block2_11 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 146:72]
        block2_11 <= block2_after_write;
      end else begin
        block2_11 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 61:26]
      block2_12 <= 512'h0; // @[DCache.scala 61:26]
    end else if (5'hc == index_addr) begin // @[DCache.scala 146:26]
      if (_T_22) begin // @[DCache.scala 146:32]
        block2_12 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 146:72]
        block2_12 <= block2_after_write;
      end else begin
        block2_12 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 61:26]
      block2_13 <= 512'h0; // @[DCache.scala 61:26]
    end else if (5'hd == index_addr) begin // @[DCache.scala 146:26]
      if (_T_22) begin // @[DCache.scala 146:32]
        block2_13 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 146:72]
        block2_13 <= block2_after_write;
      end else begin
        block2_13 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 61:26]
      block2_14 <= 512'h0; // @[DCache.scala 61:26]
    end else if (5'he == index_addr) begin // @[DCache.scala 146:26]
      if (_T_22) begin // @[DCache.scala 146:32]
        block2_14 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 146:72]
        block2_14 <= block2_after_write;
      end else begin
        block2_14 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 61:26]
      block2_15 <= 512'h0; // @[DCache.scala 61:26]
    end else if (5'hf == index_addr) begin // @[DCache.scala 146:26]
      if (_T_22) begin // @[DCache.scala 146:32]
        block2_15 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 146:72]
        block2_15 <= block2_after_write;
      end else begin
        block2_15 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 61:26]
      block2_16 <= 512'h0; // @[DCache.scala 61:26]
    end else if (5'h10 == index_addr) begin // @[DCache.scala 146:26]
      if (_T_22) begin // @[DCache.scala 146:32]
        block2_16 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 146:72]
        block2_16 <= block2_after_write;
      end else begin
        block2_16 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 61:26]
      block2_17 <= 512'h0; // @[DCache.scala 61:26]
    end else if (5'h11 == index_addr) begin // @[DCache.scala 146:26]
      if (_T_22) begin // @[DCache.scala 146:32]
        block2_17 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 146:72]
        block2_17 <= block2_after_write;
      end else begin
        block2_17 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 61:26]
      block2_18 <= 512'h0; // @[DCache.scala 61:26]
    end else if (5'h12 == index_addr) begin // @[DCache.scala 146:26]
      if (_T_22) begin // @[DCache.scala 146:32]
        block2_18 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 146:72]
        block2_18 <= block2_after_write;
      end else begin
        block2_18 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 61:26]
      block2_19 <= 512'h0; // @[DCache.scala 61:26]
    end else if (5'h13 == index_addr) begin // @[DCache.scala 146:26]
      if (_T_22) begin // @[DCache.scala 146:32]
        block2_19 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 146:72]
        block2_19 <= block2_after_write;
      end else begin
        block2_19 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 61:26]
      block2_20 <= 512'h0; // @[DCache.scala 61:26]
    end else if (5'h14 == index_addr) begin // @[DCache.scala 146:26]
      if (_T_22) begin // @[DCache.scala 146:32]
        block2_20 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 146:72]
        block2_20 <= block2_after_write;
      end else begin
        block2_20 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 61:26]
      block2_21 <= 512'h0; // @[DCache.scala 61:26]
    end else if (5'h15 == index_addr) begin // @[DCache.scala 146:26]
      if (_T_22) begin // @[DCache.scala 146:32]
        block2_21 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 146:72]
        block2_21 <= block2_after_write;
      end else begin
        block2_21 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 61:26]
      block2_22 <= 512'h0; // @[DCache.scala 61:26]
    end else if (5'h16 == index_addr) begin // @[DCache.scala 146:26]
      if (_T_22) begin // @[DCache.scala 146:32]
        block2_22 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 146:72]
        block2_22 <= block2_after_write;
      end else begin
        block2_22 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 61:26]
      block2_23 <= 512'h0; // @[DCache.scala 61:26]
    end else if (5'h17 == index_addr) begin // @[DCache.scala 146:26]
      if (_T_22) begin // @[DCache.scala 146:32]
        block2_23 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 146:72]
        block2_23 <= block2_after_write;
      end else begin
        block2_23 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 61:26]
      block2_24 <= 512'h0; // @[DCache.scala 61:26]
    end else if (5'h18 == index_addr) begin // @[DCache.scala 146:26]
      if (_T_22) begin // @[DCache.scala 146:32]
        block2_24 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 146:72]
        block2_24 <= block2_after_write;
      end else begin
        block2_24 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 61:26]
      block2_25 <= 512'h0; // @[DCache.scala 61:26]
    end else if (5'h19 == index_addr) begin // @[DCache.scala 146:26]
      if (_T_22) begin // @[DCache.scala 146:32]
        block2_25 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 146:72]
        block2_25 <= block2_after_write;
      end else begin
        block2_25 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 61:26]
      block2_26 <= 512'h0; // @[DCache.scala 61:26]
    end else if (5'h1a == index_addr) begin // @[DCache.scala 146:26]
      if (_T_22) begin // @[DCache.scala 146:32]
        block2_26 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 146:72]
        block2_26 <= block2_after_write;
      end else begin
        block2_26 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 61:26]
      block2_27 <= 512'h0; // @[DCache.scala 61:26]
    end else if (5'h1b == index_addr) begin // @[DCache.scala 146:26]
      if (_T_22) begin // @[DCache.scala 146:32]
        block2_27 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 146:72]
        block2_27 <= block2_after_write;
      end else begin
        block2_27 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 61:26]
      block2_28 <= 512'h0; // @[DCache.scala 61:26]
    end else if (5'h1c == index_addr) begin // @[DCache.scala 146:26]
      if (_T_22) begin // @[DCache.scala 146:32]
        block2_28 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 146:72]
        block2_28 <= block2_after_write;
      end else begin
        block2_28 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 61:26]
      block2_29 <= 512'h0; // @[DCache.scala 61:26]
    end else if (5'h1d == index_addr) begin // @[DCache.scala 146:26]
      if (_T_22) begin // @[DCache.scala 146:32]
        block2_29 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 146:72]
        block2_29 <= block2_after_write;
      end else begin
        block2_29 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 61:26]
      block2_30 <= 512'h0; // @[DCache.scala 61:26]
    end else if (5'h1e == index_addr) begin // @[DCache.scala 146:26]
      if (_T_22) begin // @[DCache.scala 146:32]
        block2_30 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 146:72]
        block2_30 <= block2_after_write;
      end else begin
        block2_30 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 61:26]
      block2_31 <= 512'h0; // @[DCache.scala 61:26]
    end else if (5'h1f == index_addr) begin // @[DCache.scala 146:26]
      if (_T_22) begin // @[DCache.scala 146:32]
        block2_31 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 146:72]
        block2_31 <= block2_after_write;
      end else begin
        block2_31 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 69:24]
      state <= 3'h0; // @[DCache.scala 69:24]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_fence_req) begin // @[DCache.scala 94:31]
        state <= 3'h3; // @[DCache.scala 94:38]
      end else if (miss & ~not_en_yet) begin // @[DCache.scala 95:43]
        state <= _state_T; // @[DCache.scala 95:50]
      end
    end else if (_T_3) begin // @[Conditional.scala 39:67]
      if (io_axi_wdone) begin // @[DCache.scala 98:32]
        state <= 3'h2; // @[DCache.scala 98:39]
      end
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      state <= _GEN_391;
    end else begin
      state <= _GEN_463;
    end
    not_en_yet <= reset | _not_en_yet_T; // @[DCache.scala 74:30 DCache.scala 74:30 DCache.scala 75:21]
    if (reset) begin // @[DCache.scala 91:28]
      fence_cnt <= 5'h0; // @[DCache.scala 91:28]
    end else if (_T_19 | _T_21) begin // @[DCache.scala 180:63]
      fence_cnt <= _lo_T_1; // @[DCache.scala 180:74]
    end else if (!(_T_23 | _T_25)) begin // @[DCache.scala 181:64]
      fence_cnt <= 5'h0; // @[DCache.scala 182:26]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  op = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  addr = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  wdata = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  wm = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  v1_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  v1_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  v1_2 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  v1_3 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  v1_4 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  v1_5 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  v1_6 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  v1_7 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  v1_8 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  v1_9 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  v1_10 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  v1_11 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  v1_12 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  v1_13 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  v1_14 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  v1_15 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  v1_16 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  v1_17 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  v1_18 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  v1_19 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  v1_20 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  v1_21 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  v1_22 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  v1_23 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  v1_24 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  v1_25 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  v1_26 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  v1_27 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  v1_28 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  v1_29 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  v1_30 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  v1_31 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  d1_0 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  d1_1 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  d1_2 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  d1_3 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  d1_4 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  d1_5 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  d1_6 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  d1_7 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  d1_8 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  d1_9 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  d1_10 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  d1_11 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  d1_12 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  d1_13 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  d1_14 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  d1_15 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  d1_16 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  d1_17 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  d1_18 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  d1_19 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  d1_20 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  d1_21 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  d1_22 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  d1_23 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  d1_24 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  d1_25 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  d1_26 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  d1_27 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  d1_28 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  d1_29 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  d1_30 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  d1_31 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  age1_0 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  age1_1 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  age1_2 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  age1_3 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  age1_4 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  age1_5 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  age1_6 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  age1_7 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  age1_8 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  age1_9 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  age1_10 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  age1_11 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  age1_12 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  age1_13 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  age1_14 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  age1_15 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  age1_16 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  age1_17 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  age1_18 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  age1_19 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  age1_20 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  age1_21 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  age1_22 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  age1_23 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  age1_24 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  age1_25 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  age1_26 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  age1_27 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  age1_28 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  age1_29 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  age1_30 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  age1_31 = _RAND_99[0:0];
  _RAND_100 = {2{`RANDOM}};
  tag1_0 = _RAND_100[52:0];
  _RAND_101 = {2{`RANDOM}};
  tag1_1 = _RAND_101[52:0];
  _RAND_102 = {2{`RANDOM}};
  tag1_2 = _RAND_102[52:0];
  _RAND_103 = {2{`RANDOM}};
  tag1_3 = _RAND_103[52:0];
  _RAND_104 = {2{`RANDOM}};
  tag1_4 = _RAND_104[52:0];
  _RAND_105 = {2{`RANDOM}};
  tag1_5 = _RAND_105[52:0];
  _RAND_106 = {2{`RANDOM}};
  tag1_6 = _RAND_106[52:0];
  _RAND_107 = {2{`RANDOM}};
  tag1_7 = _RAND_107[52:0];
  _RAND_108 = {2{`RANDOM}};
  tag1_8 = _RAND_108[52:0];
  _RAND_109 = {2{`RANDOM}};
  tag1_9 = _RAND_109[52:0];
  _RAND_110 = {2{`RANDOM}};
  tag1_10 = _RAND_110[52:0];
  _RAND_111 = {2{`RANDOM}};
  tag1_11 = _RAND_111[52:0];
  _RAND_112 = {2{`RANDOM}};
  tag1_12 = _RAND_112[52:0];
  _RAND_113 = {2{`RANDOM}};
  tag1_13 = _RAND_113[52:0];
  _RAND_114 = {2{`RANDOM}};
  tag1_14 = _RAND_114[52:0];
  _RAND_115 = {2{`RANDOM}};
  tag1_15 = _RAND_115[52:0];
  _RAND_116 = {2{`RANDOM}};
  tag1_16 = _RAND_116[52:0];
  _RAND_117 = {2{`RANDOM}};
  tag1_17 = _RAND_117[52:0];
  _RAND_118 = {2{`RANDOM}};
  tag1_18 = _RAND_118[52:0];
  _RAND_119 = {2{`RANDOM}};
  tag1_19 = _RAND_119[52:0];
  _RAND_120 = {2{`RANDOM}};
  tag1_20 = _RAND_120[52:0];
  _RAND_121 = {2{`RANDOM}};
  tag1_21 = _RAND_121[52:0];
  _RAND_122 = {2{`RANDOM}};
  tag1_22 = _RAND_122[52:0];
  _RAND_123 = {2{`RANDOM}};
  tag1_23 = _RAND_123[52:0];
  _RAND_124 = {2{`RANDOM}};
  tag1_24 = _RAND_124[52:0];
  _RAND_125 = {2{`RANDOM}};
  tag1_25 = _RAND_125[52:0];
  _RAND_126 = {2{`RANDOM}};
  tag1_26 = _RAND_126[52:0];
  _RAND_127 = {2{`RANDOM}};
  tag1_27 = _RAND_127[52:0];
  _RAND_128 = {2{`RANDOM}};
  tag1_28 = _RAND_128[52:0];
  _RAND_129 = {2{`RANDOM}};
  tag1_29 = _RAND_129[52:0];
  _RAND_130 = {2{`RANDOM}};
  tag1_30 = _RAND_130[52:0];
  _RAND_131 = {2{`RANDOM}};
  tag1_31 = _RAND_131[52:0];
  _RAND_132 = {16{`RANDOM}};
  block1_0 = _RAND_132[511:0];
  _RAND_133 = {16{`RANDOM}};
  block1_1 = _RAND_133[511:0];
  _RAND_134 = {16{`RANDOM}};
  block1_2 = _RAND_134[511:0];
  _RAND_135 = {16{`RANDOM}};
  block1_3 = _RAND_135[511:0];
  _RAND_136 = {16{`RANDOM}};
  block1_4 = _RAND_136[511:0];
  _RAND_137 = {16{`RANDOM}};
  block1_5 = _RAND_137[511:0];
  _RAND_138 = {16{`RANDOM}};
  block1_6 = _RAND_138[511:0];
  _RAND_139 = {16{`RANDOM}};
  block1_7 = _RAND_139[511:0];
  _RAND_140 = {16{`RANDOM}};
  block1_8 = _RAND_140[511:0];
  _RAND_141 = {16{`RANDOM}};
  block1_9 = _RAND_141[511:0];
  _RAND_142 = {16{`RANDOM}};
  block1_10 = _RAND_142[511:0];
  _RAND_143 = {16{`RANDOM}};
  block1_11 = _RAND_143[511:0];
  _RAND_144 = {16{`RANDOM}};
  block1_12 = _RAND_144[511:0];
  _RAND_145 = {16{`RANDOM}};
  block1_13 = _RAND_145[511:0];
  _RAND_146 = {16{`RANDOM}};
  block1_14 = _RAND_146[511:0];
  _RAND_147 = {16{`RANDOM}};
  block1_15 = _RAND_147[511:0];
  _RAND_148 = {16{`RANDOM}};
  block1_16 = _RAND_148[511:0];
  _RAND_149 = {16{`RANDOM}};
  block1_17 = _RAND_149[511:0];
  _RAND_150 = {16{`RANDOM}};
  block1_18 = _RAND_150[511:0];
  _RAND_151 = {16{`RANDOM}};
  block1_19 = _RAND_151[511:0];
  _RAND_152 = {16{`RANDOM}};
  block1_20 = _RAND_152[511:0];
  _RAND_153 = {16{`RANDOM}};
  block1_21 = _RAND_153[511:0];
  _RAND_154 = {16{`RANDOM}};
  block1_22 = _RAND_154[511:0];
  _RAND_155 = {16{`RANDOM}};
  block1_23 = _RAND_155[511:0];
  _RAND_156 = {16{`RANDOM}};
  block1_24 = _RAND_156[511:0];
  _RAND_157 = {16{`RANDOM}};
  block1_25 = _RAND_157[511:0];
  _RAND_158 = {16{`RANDOM}};
  block1_26 = _RAND_158[511:0];
  _RAND_159 = {16{`RANDOM}};
  block1_27 = _RAND_159[511:0];
  _RAND_160 = {16{`RANDOM}};
  block1_28 = _RAND_160[511:0];
  _RAND_161 = {16{`RANDOM}};
  block1_29 = _RAND_161[511:0];
  _RAND_162 = {16{`RANDOM}};
  block1_30 = _RAND_162[511:0];
  _RAND_163 = {16{`RANDOM}};
  block1_31 = _RAND_163[511:0];
  _RAND_164 = {1{`RANDOM}};
  v2_0 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  v2_1 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  v2_2 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  v2_3 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  v2_4 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  v2_5 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  v2_6 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  v2_7 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  v2_8 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  v2_9 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  v2_10 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  v2_11 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  v2_12 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  v2_13 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  v2_14 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  v2_15 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  v2_16 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  v2_17 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  v2_18 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  v2_19 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  v2_20 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  v2_21 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  v2_22 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  v2_23 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  v2_24 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  v2_25 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  v2_26 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  v2_27 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  v2_28 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  v2_29 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  v2_30 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  v2_31 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  d2_0 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  d2_1 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  d2_2 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  d2_3 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  d2_4 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  d2_5 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  d2_6 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  d2_7 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  d2_8 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  d2_9 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  d2_10 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  d2_11 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  d2_12 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  d2_13 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  d2_14 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  d2_15 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  d2_16 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  d2_17 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  d2_18 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  d2_19 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  d2_20 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  d2_21 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  d2_22 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  d2_23 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  d2_24 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  d2_25 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  d2_26 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  d2_27 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  d2_28 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  d2_29 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  d2_30 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  d2_31 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  age2_0 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  age2_1 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  age2_2 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  age2_3 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  age2_4 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  age2_5 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  age2_6 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  age2_7 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  age2_8 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  age2_9 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  age2_10 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  age2_11 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  age2_12 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  age2_13 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  age2_14 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  age2_15 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  age2_16 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  age2_17 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  age2_18 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  age2_19 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  age2_20 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  age2_21 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  age2_22 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  age2_23 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  age2_24 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  age2_25 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  age2_26 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  age2_27 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  age2_28 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  age2_29 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  age2_30 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  age2_31 = _RAND_259[0:0];
  _RAND_260 = {2{`RANDOM}};
  tag2_0 = _RAND_260[52:0];
  _RAND_261 = {2{`RANDOM}};
  tag2_1 = _RAND_261[52:0];
  _RAND_262 = {2{`RANDOM}};
  tag2_2 = _RAND_262[52:0];
  _RAND_263 = {2{`RANDOM}};
  tag2_3 = _RAND_263[52:0];
  _RAND_264 = {2{`RANDOM}};
  tag2_4 = _RAND_264[52:0];
  _RAND_265 = {2{`RANDOM}};
  tag2_5 = _RAND_265[52:0];
  _RAND_266 = {2{`RANDOM}};
  tag2_6 = _RAND_266[52:0];
  _RAND_267 = {2{`RANDOM}};
  tag2_7 = _RAND_267[52:0];
  _RAND_268 = {2{`RANDOM}};
  tag2_8 = _RAND_268[52:0];
  _RAND_269 = {2{`RANDOM}};
  tag2_9 = _RAND_269[52:0];
  _RAND_270 = {2{`RANDOM}};
  tag2_10 = _RAND_270[52:0];
  _RAND_271 = {2{`RANDOM}};
  tag2_11 = _RAND_271[52:0];
  _RAND_272 = {2{`RANDOM}};
  tag2_12 = _RAND_272[52:0];
  _RAND_273 = {2{`RANDOM}};
  tag2_13 = _RAND_273[52:0];
  _RAND_274 = {2{`RANDOM}};
  tag2_14 = _RAND_274[52:0];
  _RAND_275 = {2{`RANDOM}};
  tag2_15 = _RAND_275[52:0];
  _RAND_276 = {2{`RANDOM}};
  tag2_16 = _RAND_276[52:0];
  _RAND_277 = {2{`RANDOM}};
  tag2_17 = _RAND_277[52:0];
  _RAND_278 = {2{`RANDOM}};
  tag2_18 = _RAND_278[52:0];
  _RAND_279 = {2{`RANDOM}};
  tag2_19 = _RAND_279[52:0];
  _RAND_280 = {2{`RANDOM}};
  tag2_20 = _RAND_280[52:0];
  _RAND_281 = {2{`RANDOM}};
  tag2_21 = _RAND_281[52:0];
  _RAND_282 = {2{`RANDOM}};
  tag2_22 = _RAND_282[52:0];
  _RAND_283 = {2{`RANDOM}};
  tag2_23 = _RAND_283[52:0];
  _RAND_284 = {2{`RANDOM}};
  tag2_24 = _RAND_284[52:0];
  _RAND_285 = {2{`RANDOM}};
  tag2_25 = _RAND_285[52:0];
  _RAND_286 = {2{`RANDOM}};
  tag2_26 = _RAND_286[52:0];
  _RAND_287 = {2{`RANDOM}};
  tag2_27 = _RAND_287[52:0];
  _RAND_288 = {2{`RANDOM}};
  tag2_28 = _RAND_288[52:0];
  _RAND_289 = {2{`RANDOM}};
  tag2_29 = _RAND_289[52:0];
  _RAND_290 = {2{`RANDOM}};
  tag2_30 = _RAND_290[52:0];
  _RAND_291 = {2{`RANDOM}};
  tag2_31 = _RAND_291[52:0];
  _RAND_292 = {16{`RANDOM}};
  block2_0 = _RAND_292[511:0];
  _RAND_293 = {16{`RANDOM}};
  block2_1 = _RAND_293[511:0];
  _RAND_294 = {16{`RANDOM}};
  block2_2 = _RAND_294[511:0];
  _RAND_295 = {16{`RANDOM}};
  block2_3 = _RAND_295[511:0];
  _RAND_296 = {16{`RANDOM}};
  block2_4 = _RAND_296[511:0];
  _RAND_297 = {16{`RANDOM}};
  block2_5 = _RAND_297[511:0];
  _RAND_298 = {16{`RANDOM}};
  block2_6 = _RAND_298[511:0];
  _RAND_299 = {16{`RANDOM}};
  block2_7 = _RAND_299[511:0];
  _RAND_300 = {16{`RANDOM}};
  block2_8 = _RAND_300[511:0];
  _RAND_301 = {16{`RANDOM}};
  block2_9 = _RAND_301[511:0];
  _RAND_302 = {16{`RANDOM}};
  block2_10 = _RAND_302[511:0];
  _RAND_303 = {16{`RANDOM}};
  block2_11 = _RAND_303[511:0];
  _RAND_304 = {16{`RANDOM}};
  block2_12 = _RAND_304[511:0];
  _RAND_305 = {16{`RANDOM}};
  block2_13 = _RAND_305[511:0];
  _RAND_306 = {16{`RANDOM}};
  block2_14 = _RAND_306[511:0];
  _RAND_307 = {16{`RANDOM}};
  block2_15 = _RAND_307[511:0];
  _RAND_308 = {16{`RANDOM}};
  block2_16 = _RAND_308[511:0];
  _RAND_309 = {16{`RANDOM}};
  block2_17 = _RAND_309[511:0];
  _RAND_310 = {16{`RANDOM}};
  block2_18 = _RAND_310[511:0];
  _RAND_311 = {16{`RANDOM}};
  block2_19 = _RAND_311[511:0];
  _RAND_312 = {16{`RANDOM}};
  block2_20 = _RAND_312[511:0];
  _RAND_313 = {16{`RANDOM}};
  block2_21 = _RAND_313[511:0];
  _RAND_314 = {16{`RANDOM}};
  block2_22 = _RAND_314[511:0];
  _RAND_315 = {16{`RANDOM}};
  block2_23 = _RAND_315[511:0];
  _RAND_316 = {16{`RANDOM}};
  block2_24 = _RAND_316[511:0];
  _RAND_317 = {16{`RANDOM}};
  block2_25 = _RAND_317[511:0];
  _RAND_318 = {16{`RANDOM}};
  block2_26 = _RAND_318[511:0];
  _RAND_319 = {16{`RANDOM}};
  block2_27 = _RAND_319[511:0];
  _RAND_320 = {16{`RANDOM}};
  block2_28 = _RAND_320[511:0];
  _RAND_321 = {16{`RANDOM}};
  block2_29 = _RAND_321[511:0];
  _RAND_322 = {16{`RANDOM}};
  block2_30 = _RAND_322[511:0];
  _RAND_323 = {16{`RANDOM}};
  block2_31 = _RAND_323[511:0];
  _RAND_324 = {1{`RANDOM}};
  state = _RAND_324[2:0];
  _RAND_325 = {1{`RANDOM}};
  not_en_yet = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  fence_cnt = _RAND_326[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI(
  input          clock,
  input          reset,
  input          io_out_aw_ready,
  output         io_out_aw_valid,
  output [7:0]   io_out_aw_bits_len,
  output [2:0]   io_out_aw_bits_size,
  output [63:0]  io_out_aw_bits_addr,
  input          io_out_w_ready,
  output         io_out_w_valid,
  output [63:0]  io_out_w_bits_data,
  output [7:0]   io_out_w_bits_strb,
  output         io_out_w_bits_last,
  output         io_out_b_ready,
  input          io_out_b_valid,
  input          io_out_ar_ready,
  output         io_out_ar_valid,
  output [7:0]   io_out_ar_bits_len,
  output [2:0]   io_out_ar_bits_size,
  output [63:0]  io_out_ar_bits_addr,
  output         io_out_r_ready,
  input          io_out_r_valid,
  input  [63:0]  io_out_r_bits_data,
  input          io_out_r_bits_last,
  input          io_icacheio_req,
  input  [63:0]  io_icacheio_addr,
  output         io_icacheio_valid,
  output [511:0] io_icacheio_data,
  input          io_dcacheio_req,
  input  [63:0]  io_dcacheio_raddr,
  output         io_dcacheio_rvalid,
  output [511:0] io_dcacheio_rdata,
  input          io_dcacheio_weq,
  input  [63:0]  io_dcacheio_waddr,
  input  [511:0] io_dcacheio_wdata,
  output         io_dcacheio_wdone,
  input          io_icacheBypassIO_req,
  input  [31:0]  io_icacheBypassIO_addr,
  output         io_icacheBypassIO_valid,
  output [63:0]  io_icacheBypassIO_data,
  input          io_dcacheBypassIO_req,
  input  [31:0]  io_dcacheBypassIO_raddr,
  output         io_dcacheBypassIO_rvalid,
  output [63:0]  io_dcacheBypassIO_rdata,
  input          io_dcacheBypassIO_weq,
  input  [31:0]  io_dcacheBypassIO_waddr,
  input  [63:0]  io_dcacheBypassIO_wdata,
  input  [7:0]   io_dcacheBypassIO_wmask,
  output         io_dcacheBypassIO_wdone,
  input  [2:0]   io_dcacheBypassIO_transfer
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ibuffer_0; // @[AXI.scala 107:30]
  reg [63:0] ibuffer_1; // @[AXI.scala 107:30]
  reg [63:0] ibuffer_2; // @[AXI.scala 107:30]
  reg [63:0] ibuffer_3; // @[AXI.scala 107:30]
  reg [63:0] ibuffer_4; // @[AXI.scala 107:30]
  reg [63:0] ibuffer_5; // @[AXI.scala 107:30]
  reg [63:0] ibuffer_6; // @[AXI.scala 107:30]
  reg [63:0] ibuffer_7; // @[AXI.scala 107:30]
  reg [63:0] drbuffer_0; // @[AXI.scala 108:30]
  reg [63:0] drbuffer_1; // @[AXI.scala 108:30]
  reg [63:0] drbuffer_2; // @[AXI.scala 108:30]
  reg [63:0] drbuffer_3; // @[AXI.scala 108:30]
  reg [63:0] drbuffer_4; // @[AXI.scala 108:30]
  reg [63:0] drbuffer_5; // @[AXI.scala 108:30]
  reg [63:0] drbuffer_6; // @[AXI.scala 108:30]
  reg [63:0] drbuffer_7; // @[AXI.scala 108:30]
  reg [5:0] icnt; // @[AXI.scala 109:30]
  reg [5:0] drcnt; // @[AXI.scala 110:30]
  reg [5:0] dwcnt; // @[AXI.scala 111:30]
  reg [3:0] rstate; // @[AXI.scala 115:25]
  reg [2:0] wstate; // @[AXI.scala 116:25]
  reg  r_bypass; // @[AXI.scala 117:27]
  reg  w_bypass; // @[AXI.scala 118:27]
  wire  _T = 4'h0 == rstate; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_0 = io_dcacheBypassIO_req ? 4'h5 : rstate; // @[AXI.scala 135:42 AXI.scala 136:24 AXI.scala 115:25]
  wire  _GEN_1 = io_dcacheBypassIO_req | r_bypass; // @[AXI.scala 135:42 AXI.scala 137:26 AXI.scala 117:27]
  wire [3:0] _GEN_2 = io_icacheBypassIO_req ? 4'h1 : _GEN_0; // @[AXI.scala 131:42 AXI.scala 132:24]
  wire  _GEN_3 = io_icacheBypassIO_req | _GEN_1; // @[AXI.scala 131:42 AXI.scala 133:26]
  wire  _T_1 = 4'h1 == rstate; // @[Conditional.scala 37:30]
  wire  _T_2 = 4'h2 == rstate; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_9 = io_out_r_valid ? 4'h3 : rstate; // @[AXI.scala 145:31 AXI.scala 145:39 AXI.scala 115:25]
  wire  _T_3 = 4'h3 == rstate; // @[Conditional.scala 37:30]
  wire  _T_4 = io_out_r_valid & io_out_r_bits_last; // @[AXI.scala 148:30]
  wire [3:0] _GEN_10 = io_out_r_valid & io_out_r_bits_last ? 4'h4 : rstate; // @[AXI.scala 148:50 AXI.scala 148:58 AXI.scala 115:25]
  wire  _T_5 = 4'h4 == rstate; // @[Conditional.scala 37:30]
  wire  _T_6 = 4'h5 == rstate; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_11 = io_out_ar_ready ? 4'h6 : rstate; // @[AXI.scala 155:32 AXI.scala 155:40 AXI.scala 115:25]
  wire  _T_7 = 4'h6 == rstate; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_12 = io_out_r_valid ? 4'h7 : rstate; // @[AXI.scala 158:31 AXI.scala 158:39 AXI.scala 115:25]
  wire  _T_8 = 4'h7 == rstate; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_13 = _T_4 ? 4'h8 : rstate; // @[AXI.scala 161:50 AXI.scala 161:58 AXI.scala 115:25]
  wire  _T_10 = 4'h8 == rstate; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_14 = _T_10 ? 4'h0 : rstate; // @[Conditional.scala 39:67 AXI.scala 164:20 AXI.scala 115:25]
  wire [3:0] _GEN_15 = _T_8 ? _GEN_13 : _GEN_14; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_16 = _T_7 ? _GEN_12 : _GEN_15; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_17 = _T_6 ? _GEN_11 : _GEN_16; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_18 = _T_5 ? 4'h0 : _GEN_17; // @[Conditional.scala 39:67 AXI.scala 151:20]
  wire [3:0] _GEN_19 = _T_3 ? _GEN_10 : _GEN_18; // @[Conditional.scala 39:67]
  wire  _T_11 = 3'h0 == wstate; // @[Conditional.scala 37:30]
  wire  _GEN_25 = io_dcacheBypassIO_weq | w_bypass; // @[AXI.scala 175:42 AXI.scala 177:26 AXI.scala 118:27]
  wire  _T_12 = 3'h1 == wstate; // @[Conditional.scala 37:30]
  wire  _T_13 = 3'h2 == wstate; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_29 = io_out_w_bits_last & io_out_w_ready ? 3'h3 : wstate; // @[AXI.scala 184:50 AXI.scala 184:58 AXI.scala 116:25]
  wire  _T_15 = 3'h3 == wstate; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_30 = io_out_b_valid ? 3'h4 : wstate; // @[AXI.scala 187:31 AXI.scala 187:39 AXI.scala 116:25]
  wire  _T_16 = 3'h4 == wstate; // @[Conditional.scala 37:30]
  wire  _T_17 = ~io_out_b_valid; // @[AXI.scala 190:18]
  wire [2:0] _GEN_31 = ~io_out_b_valid ? 3'h0 : wstate; // @[AXI.scala 190:32 AXI.scala 190:40 AXI.scala 116:25]
  wire [2:0] _GEN_32 = _T_16 ? _GEN_31 : wstate; // @[Conditional.scala 39:67 AXI.scala 116:25]
  wire [2:0] _GEN_33 = _T_15 ? _GEN_30 : _GEN_32; // @[Conditional.scala 39:67]
  wire  _ibuffer_T = rstate == 4'h3; // @[AXI.scala 196:33]
  wire [63:0] _GEN_39 = 3'h1 == icnt[2:0] ? ibuffer_1 : ibuffer_0; // @[AXI.scala 196:25 AXI.scala 196:25]
  wire [63:0] _GEN_40 = 3'h2 == icnt[2:0] ? ibuffer_2 : _GEN_39; // @[AXI.scala 196:25 AXI.scala 196:25]
  wire [63:0] _GEN_41 = 3'h3 == icnt[2:0] ? ibuffer_3 : _GEN_40; // @[AXI.scala 196:25 AXI.scala 196:25]
  wire [63:0] _GEN_42 = 3'h4 == icnt[2:0] ? ibuffer_4 : _GEN_41; // @[AXI.scala 196:25 AXI.scala 196:25]
  wire [63:0] _GEN_43 = 3'h5 == icnt[2:0] ? ibuffer_5 : _GEN_42; // @[AXI.scala 196:25 AXI.scala 196:25]
  wire [63:0] _GEN_44 = 3'h6 == icnt[2:0] ? ibuffer_6 : _GEN_43; // @[AXI.scala 196:25 AXI.scala 196:25]
  wire [5:0] _icnt_T_2 = icnt + 6'h1; // @[AXI.scala 197:59]
  wire  _drbuffer_T = rstate == 4'h7; // @[AXI.scala 198:35]
  wire [63:0] _GEN_55 = 3'h1 == drcnt[2:0] ? drbuffer_1 : drbuffer_0; // @[AXI.scala 198:27 AXI.scala 198:27]
  wire [63:0] _GEN_56 = 3'h2 == drcnt[2:0] ? drbuffer_2 : _GEN_55; // @[AXI.scala 198:27 AXI.scala 198:27]
  wire [63:0] _GEN_57 = 3'h3 == drcnt[2:0] ? drbuffer_3 : _GEN_56; // @[AXI.scala 198:27 AXI.scala 198:27]
  wire [63:0] _GEN_58 = 3'h4 == drcnt[2:0] ? drbuffer_4 : _GEN_57; // @[AXI.scala 198:27 AXI.scala 198:27]
  wire [63:0] _GEN_59 = 3'h5 == drcnt[2:0] ? drbuffer_5 : _GEN_58; // @[AXI.scala 198:27 AXI.scala 198:27]
  wire [63:0] _GEN_60 = 3'h6 == drcnt[2:0] ? drbuffer_6 : _GEN_59; // @[AXI.scala 198:27 AXI.scala 198:27]
  wire [5:0] _drcnt_T_2 = drcnt + 6'h1; // @[AXI.scala 199:61]
  wire [5:0] _dwcnt_T_2 = dwcnt + 6'h1; // @[AXI.scala 200:60]
  wire [512:0] _T_20 = {ibuffer_7,ibuffer_6,ibuffer_5,ibuffer_4,ibuffer_3,ibuffer_2,ibuffer_1,ibuffer_0,1'h0}; // @[Cat.scala 30:58]
  wire [511:0] idata = _T_20[512:1]; // @[AXI.scala 206:18]
  wire [512:0] _T_21 = {drbuffer_7,drbuffer_6,drbuffer_5,drbuffer_4,drbuffer_3,drbuffer_2,drbuffer_1,drbuffer_0,1'h0}; // @[Cat.scala 30:58]
  wire [511:0] drdata = _T_21[512:1]; // @[AXI.scala 209:20]
  wire  _io_icacheio_valid_T = rstate == 4'h4; // @[AXI.scala 214:31]
  wire  _io_icacheio_valid_T_1 = ~r_bypass; // @[AXI.scala 214:55]
  wire  _io_dcacheio_rvalid_T = rstate == 4'h8; // @[AXI.scala 219:31]
  wire  _io_dcacheio_wdone_T_2 = wstate == 3'h4 & _T_17; // @[AXI.scala 221:42]
  wire  sel_raddr_hi_hi = rstate == 4'h1; // @[AXI.scala 237:32]
  wire  sel_raddr_hi_lo = rstate == 4'h5; // @[AXI.scala 237:52]
  wire [2:0] sel_raddr = {sel_raddr_hi_hi,sel_raddr_hi_lo,r_bypass}; // @[Cat.scala 30:58]
  wire [63:0] _io_out_ar_bits_addr_T_1 = 3'h4 == sel_raddr ? io_icacheio_addr : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _io_out_ar_bits_addr_T_3 = 3'h2 == sel_raddr ? io_dcacheio_raddr : _io_out_ar_bits_addr_T_1; // @[Mux.scala 80:57]
  wire [63:0] _io_out_ar_bits_addr_T_5 = 3'h5 == sel_raddr ? {{32'd0}, io_icacheBypassIO_addr} :
    _io_out_ar_bits_addr_T_3; // @[Mux.scala 80:57]
  wire [2:0] _io_out_ar_bits_len_T = r_bypass ? 3'h0 : 3'h7; // @[AXI.scala 250:31]
  wire [1:0] _io_out_ar_bits_size_T_1 = 3'h4 == sel_raddr ? 2'h3 : 2'h0; // @[Mux.scala 80:57]
  wire [1:0] _io_out_ar_bits_size_T_3 = 3'h2 == sel_raddr ? 2'h3 : _io_out_ar_bits_size_T_1; // @[Mux.scala 80:57]
  wire [1:0] _io_out_ar_bits_size_T_5 = 3'h5 == sel_raddr ? 2'h2 : _io_out_ar_bits_size_T_3; // @[Mux.scala 80:57]
  wire [2:0] _io_out_aw_bits_len_T = w_bypass ? 3'h0 : 3'h7; // @[AXI.scala 278:31]
  wire [11:0] _io_out_w_bits_data_T = {dwcnt, 6'h0}; // @[AXI.scala 286:90]
  wire [511:0] _io_out_w_bits_data_T_1 = io_dcacheio_wdata >> _io_out_w_bits_data_T; // @[AXI.scala 286:80]
  assign io_out_aw_valid = wstate == 3'h1; // @[AXI.scala 273:35]
  assign io_out_aw_bits_len = {{5'd0}, _io_out_aw_bits_len_T}; // @[AXI.scala 278:31]
  assign io_out_aw_bits_size = w_bypass ? io_dcacheBypassIO_transfer : 3'h3; // @[AXI.scala 279:31]
  assign io_out_aw_bits_addr = w_bypass ? {{32'd0}, io_dcacheBypassIO_waddr} : io_dcacheio_waddr; // @[AXI.scala 274:31]
  assign io_out_w_valid = wstate == 3'h2; // @[AXI.scala 285:35]
  assign io_out_w_bits_data = w_bypass ? io_dcacheBypassIO_wdata : _io_out_w_bits_data_T_1[63:0]; // @[AXI.scala 286:31]
  assign io_out_w_bits_strb = w_bypass ? io_dcacheBypassIO_wmask : 8'hff; // @[AXI.scala 287:31]
  assign io_out_w_bits_last = w_bypass ? dwcnt == 6'h0 : dwcnt == 6'h7; // @[AXI.scala 288:31]
  assign io_out_b_ready = wstate == 3'h4; // @[AXI.scala 290:35]
  assign io_out_ar_valid = sel_raddr_hi_hi | sel_raddr_hi_lo; // @[AXI.scala 240:47]
  assign io_out_ar_bits_len = {{5'd0}, _io_out_ar_bits_len_T}; // @[AXI.scala 250:31]
  assign io_out_ar_bits_size = 3'h3 == sel_raddr ? io_dcacheBypassIO_transfer : {{1'd0}, _io_out_ar_bits_size_T_5}; // @[Mux.scala 80:57]
  assign io_out_ar_bits_addr = 3'h3 == sel_raddr ? {{32'd0}, io_dcacheBypassIO_raddr} : _io_out_ar_bits_addr_T_5; // @[Mux.scala 80:57]
  assign io_out_r_ready = _ibuffer_T | _drbuffer_T; // @[AXI.scala 269:47]
  assign io_icacheio_valid = rstate == 4'h4 & ~r_bypass; // @[AXI.scala 214:43]
  assign io_icacheio_data = _T_20[512:1]; // @[AXI.scala 206:18]
  assign io_dcacheio_rvalid = rstate == 4'h8 & _io_icacheio_valid_T_1; // @[AXI.scala 219:43]
  assign io_dcacheio_rdata = _T_21[512:1]; // @[AXI.scala 209:20]
  assign io_dcacheio_wdone = wstate == 3'h4 & _T_17; // @[AXI.scala 221:42]
  assign io_icacheBypassIO_valid = _io_icacheio_valid_T & r_bypass; // @[AXI.scala 225:49]
  assign io_icacheBypassIO_data = idata[63:0]; // @[AXI.scala 226:35]
  assign io_dcacheBypassIO_rvalid = _io_dcacheio_rvalid_T & r_bypass; // @[AXI.scala 231:49]
  assign io_dcacheBypassIO_rdata = drdata[63:0]; // @[AXI.scala 232:36]
  assign io_dcacheBypassIO_wdone = _io_dcacheio_wdone_T_2 & w_bypass; // @[AXI.scala 233:64]
  always @(posedge clock) begin
    if (reset) begin // @[AXI.scala 107:30]
      ibuffer_0 <= 64'h0; // @[AXI.scala 107:30]
    end else if (3'h0 == icnt[2:0]) begin // @[AXI.scala 196:19]
      if (rstate == 4'h3) begin // @[AXI.scala 196:25]
        ibuffer_0 <= io_out_r_bits_data;
      end else if (3'h7 == icnt[2:0]) begin // @[AXI.scala 196:25]
        ibuffer_0 <= ibuffer_7; // @[AXI.scala 196:25]
      end else begin
        ibuffer_0 <= _GEN_44;
      end
    end
    if (reset) begin // @[AXI.scala 107:30]
      ibuffer_1 <= 64'h0; // @[AXI.scala 107:30]
    end else if (3'h1 == icnt[2:0]) begin // @[AXI.scala 196:19]
      if (rstate == 4'h3) begin // @[AXI.scala 196:25]
        ibuffer_1 <= io_out_r_bits_data;
      end else if (3'h7 == icnt[2:0]) begin // @[AXI.scala 196:25]
        ibuffer_1 <= ibuffer_7; // @[AXI.scala 196:25]
      end else begin
        ibuffer_1 <= _GEN_44;
      end
    end
    if (reset) begin // @[AXI.scala 107:30]
      ibuffer_2 <= 64'h0; // @[AXI.scala 107:30]
    end else if (3'h2 == icnt[2:0]) begin // @[AXI.scala 196:19]
      if (rstate == 4'h3) begin // @[AXI.scala 196:25]
        ibuffer_2 <= io_out_r_bits_data;
      end else if (3'h7 == icnt[2:0]) begin // @[AXI.scala 196:25]
        ibuffer_2 <= ibuffer_7; // @[AXI.scala 196:25]
      end else begin
        ibuffer_2 <= _GEN_44;
      end
    end
    if (reset) begin // @[AXI.scala 107:30]
      ibuffer_3 <= 64'h0; // @[AXI.scala 107:30]
    end else if (3'h3 == icnt[2:0]) begin // @[AXI.scala 196:19]
      if (rstate == 4'h3) begin // @[AXI.scala 196:25]
        ibuffer_3 <= io_out_r_bits_data;
      end else if (3'h7 == icnt[2:0]) begin // @[AXI.scala 196:25]
        ibuffer_3 <= ibuffer_7; // @[AXI.scala 196:25]
      end else begin
        ibuffer_3 <= _GEN_44;
      end
    end
    if (reset) begin // @[AXI.scala 107:30]
      ibuffer_4 <= 64'h0; // @[AXI.scala 107:30]
    end else if (3'h4 == icnt[2:0]) begin // @[AXI.scala 196:19]
      if (rstate == 4'h3) begin // @[AXI.scala 196:25]
        ibuffer_4 <= io_out_r_bits_data;
      end else if (3'h7 == icnt[2:0]) begin // @[AXI.scala 196:25]
        ibuffer_4 <= ibuffer_7; // @[AXI.scala 196:25]
      end else begin
        ibuffer_4 <= _GEN_44;
      end
    end
    if (reset) begin // @[AXI.scala 107:30]
      ibuffer_5 <= 64'h0; // @[AXI.scala 107:30]
    end else if (3'h5 == icnt[2:0]) begin // @[AXI.scala 196:19]
      if (rstate == 4'h3) begin // @[AXI.scala 196:25]
        ibuffer_5 <= io_out_r_bits_data;
      end else if (3'h7 == icnt[2:0]) begin // @[AXI.scala 196:25]
        ibuffer_5 <= ibuffer_7; // @[AXI.scala 196:25]
      end else begin
        ibuffer_5 <= _GEN_44;
      end
    end
    if (reset) begin // @[AXI.scala 107:30]
      ibuffer_6 <= 64'h0; // @[AXI.scala 107:30]
    end else if (3'h6 == icnt[2:0]) begin // @[AXI.scala 196:19]
      if (rstate == 4'h3) begin // @[AXI.scala 196:25]
        ibuffer_6 <= io_out_r_bits_data;
      end else if (3'h7 == icnt[2:0]) begin // @[AXI.scala 196:25]
        ibuffer_6 <= ibuffer_7; // @[AXI.scala 196:25]
      end else begin
        ibuffer_6 <= _GEN_44;
      end
    end
    if (reset) begin // @[AXI.scala 107:30]
      ibuffer_7 <= 64'h0; // @[AXI.scala 107:30]
    end else if (3'h7 == icnt[2:0]) begin // @[AXI.scala 196:19]
      if (rstate == 4'h3) begin // @[AXI.scala 196:25]
        ibuffer_7 <= io_out_r_bits_data;
      end else if (!(3'h7 == icnt[2:0])) begin // @[AXI.scala 196:25]
        ibuffer_7 <= _GEN_44;
      end
    end
    if (reset) begin // @[AXI.scala 108:30]
      drbuffer_0 <= 64'h0; // @[AXI.scala 108:30]
    end else if (3'h0 == drcnt[2:0]) begin // @[AXI.scala 198:21]
      if (rstate == 4'h7) begin // @[AXI.scala 198:27]
        drbuffer_0 <= io_out_r_bits_data;
      end else if (3'h7 == drcnt[2:0]) begin // @[AXI.scala 198:27]
        drbuffer_0 <= drbuffer_7; // @[AXI.scala 198:27]
      end else begin
        drbuffer_0 <= _GEN_60;
      end
    end
    if (reset) begin // @[AXI.scala 108:30]
      drbuffer_1 <= 64'h0; // @[AXI.scala 108:30]
    end else if (3'h1 == drcnt[2:0]) begin // @[AXI.scala 198:21]
      if (rstate == 4'h7) begin // @[AXI.scala 198:27]
        drbuffer_1 <= io_out_r_bits_data;
      end else if (3'h7 == drcnt[2:0]) begin // @[AXI.scala 198:27]
        drbuffer_1 <= drbuffer_7; // @[AXI.scala 198:27]
      end else begin
        drbuffer_1 <= _GEN_60;
      end
    end
    if (reset) begin // @[AXI.scala 108:30]
      drbuffer_2 <= 64'h0; // @[AXI.scala 108:30]
    end else if (3'h2 == drcnt[2:0]) begin // @[AXI.scala 198:21]
      if (rstate == 4'h7) begin // @[AXI.scala 198:27]
        drbuffer_2 <= io_out_r_bits_data;
      end else if (3'h7 == drcnt[2:0]) begin // @[AXI.scala 198:27]
        drbuffer_2 <= drbuffer_7; // @[AXI.scala 198:27]
      end else begin
        drbuffer_2 <= _GEN_60;
      end
    end
    if (reset) begin // @[AXI.scala 108:30]
      drbuffer_3 <= 64'h0; // @[AXI.scala 108:30]
    end else if (3'h3 == drcnt[2:0]) begin // @[AXI.scala 198:21]
      if (rstate == 4'h7) begin // @[AXI.scala 198:27]
        drbuffer_3 <= io_out_r_bits_data;
      end else if (3'h7 == drcnt[2:0]) begin // @[AXI.scala 198:27]
        drbuffer_3 <= drbuffer_7; // @[AXI.scala 198:27]
      end else begin
        drbuffer_3 <= _GEN_60;
      end
    end
    if (reset) begin // @[AXI.scala 108:30]
      drbuffer_4 <= 64'h0; // @[AXI.scala 108:30]
    end else if (3'h4 == drcnt[2:0]) begin // @[AXI.scala 198:21]
      if (rstate == 4'h7) begin // @[AXI.scala 198:27]
        drbuffer_4 <= io_out_r_bits_data;
      end else if (3'h7 == drcnt[2:0]) begin // @[AXI.scala 198:27]
        drbuffer_4 <= drbuffer_7; // @[AXI.scala 198:27]
      end else begin
        drbuffer_4 <= _GEN_60;
      end
    end
    if (reset) begin // @[AXI.scala 108:30]
      drbuffer_5 <= 64'h0; // @[AXI.scala 108:30]
    end else if (3'h5 == drcnt[2:0]) begin // @[AXI.scala 198:21]
      if (rstate == 4'h7) begin // @[AXI.scala 198:27]
        drbuffer_5 <= io_out_r_bits_data;
      end else if (3'h7 == drcnt[2:0]) begin // @[AXI.scala 198:27]
        drbuffer_5 <= drbuffer_7; // @[AXI.scala 198:27]
      end else begin
        drbuffer_5 <= _GEN_60;
      end
    end
    if (reset) begin // @[AXI.scala 108:30]
      drbuffer_6 <= 64'h0; // @[AXI.scala 108:30]
    end else if (3'h6 == drcnt[2:0]) begin // @[AXI.scala 198:21]
      if (rstate == 4'h7) begin // @[AXI.scala 198:27]
        drbuffer_6 <= io_out_r_bits_data;
      end else if (3'h7 == drcnt[2:0]) begin // @[AXI.scala 198:27]
        drbuffer_6 <= drbuffer_7; // @[AXI.scala 198:27]
      end else begin
        drbuffer_6 <= _GEN_60;
      end
    end
    if (reset) begin // @[AXI.scala 108:30]
      drbuffer_7 <= 64'h0; // @[AXI.scala 108:30]
    end else if (3'h7 == drcnt[2:0]) begin // @[AXI.scala 198:21]
      if (rstate == 4'h7) begin // @[AXI.scala 198:27]
        drbuffer_7 <= io_out_r_bits_data;
      end else if (!(3'h7 == drcnt[2:0])) begin // @[AXI.scala 198:27]
        drbuffer_7 <= _GEN_60;
      end
    end
    if (reset) begin // @[AXI.scala 109:30]
      icnt <= 6'h0; // @[AXI.scala 109:30]
    end else if (_ibuffer_T) begin // @[AXI.scala 197:16]
      if (io_out_r_valid) begin // @[AXI.scala 197:40]
        icnt <= _icnt_T_2;
      end
    end else begin
      icnt <= 6'h0;
    end
    if (reset) begin // @[AXI.scala 110:30]
      drcnt <= 6'h0; // @[AXI.scala 110:30]
    end else if (_drbuffer_T) begin // @[AXI.scala 199:17]
      if (io_out_r_valid) begin // @[AXI.scala 199:41]
        drcnt <= _drcnt_T_2;
      end
    end else begin
      drcnt <= 6'h0;
    end
    if (reset) begin // @[AXI.scala 111:30]
      dwcnt <= 6'h0; // @[AXI.scala 111:30]
    end else if (wstate == 3'h2) begin // @[AXI.scala 200:17]
      if (io_out_w_ready) begin // @[AXI.scala 200:40]
        dwcnt <= _dwcnt_T_2;
      end
    end else begin
      dwcnt <= 6'h0;
    end
    if (reset) begin // @[AXI.scala 115:25]
      rstate <= 4'h0; // @[AXI.scala 115:25]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_icacheio_req) begin // @[AXI.scala 123:31]
        rstate <= 4'h1; // @[AXI.scala 124:24]
      end else if (io_dcacheio_req) begin // @[AXI.scala 127:36]
        rstate <= 4'h5; // @[AXI.scala 128:24]
      end else begin
        rstate <= _GEN_2;
      end
    end else if (_T_1) begin // @[Conditional.scala 39:67]
      if (io_out_ar_ready) begin // @[AXI.scala 142:32]
        rstate <= 4'h2; // @[AXI.scala 142:40]
      end
    end else if (_T_2) begin // @[Conditional.scala 39:67]
      rstate <= _GEN_9;
    end else begin
      rstate <= _GEN_19;
    end
    if (reset) begin // @[AXI.scala 116:25]
      wstate <= 3'h0; // @[AXI.scala 116:25]
    end else if (_T_11) begin // @[Conditional.scala 40:58]
      if (io_dcacheio_weq) begin // @[AXI.scala 171:31]
        wstate <= 3'h1; // @[AXI.scala 172:24]
      end else if (io_dcacheBypassIO_weq) begin // @[AXI.scala 175:42]
        wstate <= 3'h1; // @[AXI.scala 176:24]
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      if (io_out_aw_ready) begin // @[AXI.scala 181:32]
        wstate <= 3'h2; // @[AXI.scala 181:40]
      end
    end else if (_T_13) begin // @[Conditional.scala 39:67]
      wstate <= _GEN_29;
    end else begin
      wstate <= _GEN_33;
    end
    if (reset) begin // @[AXI.scala 117:27]
      r_bypass <= 1'h0; // @[AXI.scala 117:27]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_icacheio_req) begin // @[AXI.scala 123:31]
        r_bypass <= 1'h0; // @[AXI.scala 125:26]
      end else if (io_dcacheio_req) begin // @[AXI.scala 127:36]
        r_bypass <= 1'h0; // @[AXI.scala 129:26]
      end else begin
        r_bypass <= _GEN_3;
      end
    end
    if (reset) begin // @[AXI.scala 118:27]
      w_bypass <= 1'h0; // @[AXI.scala 118:27]
    end else if (_T_11) begin // @[Conditional.scala 40:58]
      if (io_dcacheio_weq) begin // @[AXI.scala 171:31]
        w_bypass <= 1'h0; // @[AXI.scala 173:26]
      end else begin
        w_bypass <= _GEN_25;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  ibuffer_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  ibuffer_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  ibuffer_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  ibuffer_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  ibuffer_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  ibuffer_5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  ibuffer_6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  ibuffer_7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  drbuffer_0 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  drbuffer_1 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  drbuffer_2 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  drbuffer_3 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  drbuffer_4 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  drbuffer_5 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  drbuffer_6 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  drbuffer_7 = _RAND_15[63:0];
  _RAND_16 = {1{`RANDOM}};
  icnt = _RAND_16[5:0];
  _RAND_17 = {1{`RANDOM}};
  drcnt = _RAND_17[5:0];
  _RAND_18 = {1{`RANDOM}};
  dwcnt = _RAND_18[5:0];
  _RAND_19 = {1{`RANDOM}};
  rstate = _RAND_19[3:0];
  _RAND_20 = {1{`RANDOM}};
  wstate = _RAND_20[2:0];
  _RAND_21 = {1{`RANDOM}};
  r_bypass = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  w_bypass = _RAND_22[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ICacheSocAxi(
  input          clock,
  input          reset,
  input          io_in_req,
  input  [63:0]  io_in_addr,
  output         io_in_valid,
  output [511:0] io_in_data,
  output         io_out0_req,
  output [63:0]  io_out0_addr,
  input          io_out0_valid,
  input  [511:0] io_out0_data,
  output         io_out1_req,
  output [31:0]  io_out1_addr,
  input          io_out1_valid,
  input  [63:0]  io_out1_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[CacheBypass.scala 131:24]
  reg [3:0] cnt; // @[CacheBypass.scala 133:22]
  reg [31:0] buffer_0; // @[CacheBypass.scala 134:25]
  reg [31:0] buffer_1; // @[CacheBypass.scala 134:25]
  reg [31:0] buffer_2; // @[CacheBypass.scala 134:25]
  reg [31:0] buffer_3; // @[CacheBypass.scala 134:25]
  reg [31:0] buffer_4; // @[CacheBypass.scala 134:25]
  reg [31:0] buffer_5; // @[CacheBypass.scala 134:25]
  reg [31:0] buffer_6; // @[CacheBypass.scala 134:25]
  reg [31:0] buffer_7; // @[CacheBypass.scala 134:25]
  reg [31:0] buffer_8; // @[CacheBypass.scala 134:25]
  reg [31:0] buffer_9; // @[CacheBypass.scala 134:25]
  reg [31:0] buffer_10; // @[CacheBypass.scala 134:25]
  reg [31:0] buffer_11; // @[CacheBypass.scala 134:25]
  reg [31:0] buffer_12; // @[CacheBypass.scala 134:25]
  reg [31:0] buffer_13; // @[CacheBypass.scala 134:25]
  reg [31:0] buffer_14; // @[CacheBypass.scala 134:25]
  reg [31:0] buffer_15; // @[CacheBypass.scala 134:25]
  wire  _T = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_3 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_4 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_5 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_3 = io_out1_valid ? 3'h4 : state; // @[CacheBypass.scala 149:32 CacheBypass.scala 149:39 CacheBypass.scala 131:24]
  wire  _T_6 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_4 = cnt == 4'hf ? 3'h5 : 3'h3; // @[CacheBypass.scala 152:40 CacheBypass.scala 152:47 CacheBypass.scala 153:30]
  wire  _T_8 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_5 = _T_8 ? 3'h0 : state; // @[Conditional.scala 39:67 CacheBypass.scala 156:19 CacheBypass.scala 131:24]
  wire [2:0] _GEN_6 = _T_6 ? _GEN_4 : _GEN_5; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_7 = _T_5 ? _GEN_3 : _GEN_6; // @[Conditional.scala 39:67]
  wire  _T_9 = state == 3'h4; // @[CacheBypass.scala 160:16]
  wire [288:0] lo_8 = {buffer_8,buffer_7,buffer_6,buffer_5,buffer_4,buffer_3,buffer_2,buffer_1,buffer_0,1'h0}; // @[Cat.scala 30:58]
  wire [512:0] _T_10 = {buffer_15,buffer_14,buffer_13,buffer_12,buffer_11,buffer_10,buffer_9,lo_8}; // @[Cat.scala 30:58]
  wire [511:0] data = _T_10[512:1]; // @[CacheBypass.scala 163:16]
  wire [3:0] _cnt_T_1 = cnt + 4'h1; // @[CacheBypass.scala 165:41]
  wire  _T_12 = state == 3'h5; // @[CacheBypass.scala 166:21]
  wire [5:0] _GEN_47 = {cnt, 2'h0}; // @[CacheBypass.scala 172:39]
  wire [6:0] _io_out1_addr_T = {{1'd0}, _GEN_47}; // @[CacheBypass.scala 172:39]
  wire [63:0] _GEN_48 = {{57'd0}, _io_out1_addr_T}; // @[CacheBypass.scala 172:32]
  wire [63:0] _io_out1_addr_T_2 = io_in_addr + _GEN_48; // @[CacheBypass.scala 172:32]
  wire  _io_in_valid_T_1 = state == 3'h2; // @[CacheBypass.scala 174:52]
  wire [511:0] _GEN_45 = _T_12 ? data : 512'h0; // @[CacheBypass.scala 176:38 CacheBypass.scala 176:50 CacheBypass.scala 177:27]
  assign io_in_valid = _T_12 | state == 3'h2; // @[CacheBypass.scala 174:43]
  assign io_in_data = _io_in_valid_T_1 ? io_out0_data : _GEN_45; // @[CacheBypass.scala 175:25 CacheBypass.scala 175:37]
  assign io_out0_req = state == 3'h1; // @[CacheBypass.scala 169:27]
  assign io_out0_addr = io_in_addr; // @[CacheBypass.scala 170:18]
  assign io_out1_req = state == 3'h3; // @[CacheBypass.scala 171:27]
  assign io_out1_addr = _io_out1_addr_T_2[31:0]; // @[CacheBypass.scala 172:18]
  always @(posedge clock) begin
    if (reset) begin // @[CacheBypass.scala 131:24]
      state <= 3'h0; // @[CacheBypass.scala 131:24]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_in_req & io_in_addr < 64'h80000000) begin // @[CacheBypass.scala 138:60]
        state <= 3'h3; // @[CacheBypass.scala 138:67]
      end else if (io_in_req) begin // @[CacheBypass.scala 139:33]
        state <= 3'h1; // @[CacheBypass.scala 139:40]
      end
    end else if (_T_3) begin // @[Conditional.scala 39:67]
      if (io_out0_valid) begin // @[CacheBypass.scala 143:32]
        state <= 3'h2; // @[CacheBypass.scala 143:39]
      end
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      state <= 3'h0; // @[CacheBypass.scala 146:19]
    end else begin
      state <= _GEN_7;
    end
    if (reset) begin // @[CacheBypass.scala 133:22]
      cnt <= 4'h0; // @[CacheBypass.scala 133:22]
    end else if (_T_9) begin // @[CacheBypass.scala 165:29]
      cnt <= _cnt_T_1; // @[CacheBypass.scala 165:34]
    end else if (state == 3'h5) begin // @[CacheBypass.scala 166:38]
      cnt <= 4'h0; // @[CacheBypass.scala 166:43]
    end
    if (reset) begin // @[CacheBypass.scala 134:25]
      buffer_0 <= 32'h0; // @[CacheBypass.scala 134:25]
    end else if (state == 3'h4) begin // @[CacheBypass.scala 160:29]
      if (4'h0 == cnt) begin // @[CacheBypass.scala 160:42]
        buffer_0 <= io_out1_data[31:0]; // @[CacheBypass.scala 160:42]
      end
    end
    if (reset) begin // @[CacheBypass.scala 134:25]
      buffer_1 <= 32'h0; // @[CacheBypass.scala 134:25]
    end else if (state == 3'h4) begin // @[CacheBypass.scala 160:29]
      if (4'h1 == cnt) begin // @[CacheBypass.scala 160:42]
        buffer_1 <= io_out1_data[31:0]; // @[CacheBypass.scala 160:42]
      end
    end
    if (reset) begin // @[CacheBypass.scala 134:25]
      buffer_2 <= 32'h0; // @[CacheBypass.scala 134:25]
    end else if (state == 3'h4) begin // @[CacheBypass.scala 160:29]
      if (4'h2 == cnt) begin // @[CacheBypass.scala 160:42]
        buffer_2 <= io_out1_data[31:0]; // @[CacheBypass.scala 160:42]
      end
    end
    if (reset) begin // @[CacheBypass.scala 134:25]
      buffer_3 <= 32'h0; // @[CacheBypass.scala 134:25]
    end else if (state == 3'h4) begin // @[CacheBypass.scala 160:29]
      if (4'h3 == cnt) begin // @[CacheBypass.scala 160:42]
        buffer_3 <= io_out1_data[31:0]; // @[CacheBypass.scala 160:42]
      end
    end
    if (reset) begin // @[CacheBypass.scala 134:25]
      buffer_4 <= 32'h0; // @[CacheBypass.scala 134:25]
    end else if (state == 3'h4) begin // @[CacheBypass.scala 160:29]
      if (4'h4 == cnt) begin // @[CacheBypass.scala 160:42]
        buffer_4 <= io_out1_data[31:0]; // @[CacheBypass.scala 160:42]
      end
    end
    if (reset) begin // @[CacheBypass.scala 134:25]
      buffer_5 <= 32'h0; // @[CacheBypass.scala 134:25]
    end else if (state == 3'h4) begin // @[CacheBypass.scala 160:29]
      if (4'h5 == cnt) begin // @[CacheBypass.scala 160:42]
        buffer_5 <= io_out1_data[31:0]; // @[CacheBypass.scala 160:42]
      end
    end
    if (reset) begin // @[CacheBypass.scala 134:25]
      buffer_6 <= 32'h0; // @[CacheBypass.scala 134:25]
    end else if (state == 3'h4) begin // @[CacheBypass.scala 160:29]
      if (4'h6 == cnt) begin // @[CacheBypass.scala 160:42]
        buffer_6 <= io_out1_data[31:0]; // @[CacheBypass.scala 160:42]
      end
    end
    if (reset) begin // @[CacheBypass.scala 134:25]
      buffer_7 <= 32'h0; // @[CacheBypass.scala 134:25]
    end else if (state == 3'h4) begin // @[CacheBypass.scala 160:29]
      if (4'h7 == cnt) begin // @[CacheBypass.scala 160:42]
        buffer_7 <= io_out1_data[31:0]; // @[CacheBypass.scala 160:42]
      end
    end
    if (reset) begin // @[CacheBypass.scala 134:25]
      buffer_8 <= 32'h0; // @[CacheBypass.scala 134:25]
    end else if (state == 3'h4) begin // @[CacheBypass.scala 160:29]
      if (4'h8 == cnt) begin // @[CacheBypass.scala 160:42]
        buffer_8 <= io_out1_data[31:0]; // @[CacheBypass.scala 160:42]
      end
    end
    if (reset) begin // @[CacheBypass.scala 134:25]
      buffer_9 <= 32'h0; // @[CacheBypass.scala 134:25]
    end else if (state == 3'h4) begin // @[CacheBypass.scala 160:29]
      if (4'h9 == cnt) begin // @[CacheBypass.scala 160:42]
        buffer_9 <= io_out1_data[31:0]; // @[CacheBypass.scala 160:42]
      end
    end
    if (reset) begin // @[CacheBypass.scala 134:25]
      buffer_10 <= 32'h0; // @[CacheBypass.scala 134:25]
    end else if (state == 3'h4) begin // @[CacheBypass.scala 160:29]
      if (4'ha == cnt) begin // @[CacheBypass.scala 160:42]
        buffer_10 <= io_out1_data[31:0]; // @[CacheBypass.scala 160:42]
      end
    end
    if (reset) begin // @[CacheBypass.scala 134:25]
      buffer_11 <= 32'h0; // @[CacheBypass.scala 134:25]
    end else if (state == 3'h4) begin // @[CacheBypass.scala 160:29]
      if (4'hb == cnt) begin // @[CacheBypass.scala 160:42]
        buffer_11 <= io_out1_data[31:0]; // @[CacheBypass.scala 160:42]
      end
    end
    if (reset) begin // @[CacheBypass.scala 134:25]
      buffer_12 <= 32'h0; // @[CacheBypass.scala 134:25]
    end else if (state == 3'h4) begin // @[CacheBypass.scala 160:29]
      if (4'hc == cnt) begin // @[CacheBypass.scala 160:42]
        buffer_12 <= io_out1_data[31:0]; // @[CacheBypass.scala 160:42]
      end
    end
    if (reset) begin // @[CacheBypass.scala 134:25]
      buffer_13 <= 32'h0; // @[CacheBypass.scala 134:25]
    end else if (state == 3'h4) begin // @[CacheBypass.scala 160:29]
      if (4'hd == cnt) begin // @[CacheBypass.scala 160:42]
        buffer_13 <= io_out1_data[31:0]; // @[CacheBypass.scala 160:42]
      end
    end
    if (reset) begin // @[CacheBypass.scala 134:25]
      buffer_14 <= 32'h0; // @[CacheBypass.scala 134:25]
    end else if (state == 3'h4) begin // @[CacheBypass.scala 160:29]
      if (4'he == cnt) begin // @[CacheBypass.scala 160:42]
        buffer_14 <= io_out1_data[31:0]; // @[CacheBypass.scala 160:42]
      end
    end
    if (reset) begin // @[CacheBypass.scala 134:25]
      buffer_15 <= 32'h0; // @[CacheBypass.scala 134:25]
    end else if (state == 3'h4) begin // @[CacheBypass.scala 160:29]
      if (4'hf == cnt) begin // @[CacheBypass.scala 160:42]
        buffer_15 <= io_out1_data[31:0]; // @[CacheBypass.scala 160:42]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  cnt = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  buffer_0 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  buffer_1 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  buffer_2 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  buffer_3 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  buffer_4 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  buffer_5 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  buffer_6 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  buffer_7 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  buffer_8 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  buffer_9 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  buffer_10 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  buffer_11 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  buffer_12 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  buffer_13 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  buffer_14 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  buffer_15 = _RAND_17[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DMMIO(
  input         clock,
  input         reset,
  input         io_dmem_en,
  input         io_dmem_op,
  input  [63:0] io_dmem_addr,
  input  [63:0] io_dmem_wdata,
  input  [7:0]  io_dmem_wmask,
  input  [31:0] io_dmem_transfer,
  output        io_dmem_ok,
  output [63:0] io_dmem_rdata,
  output        io_mem0_en,
  output        io_mem0_op,
  output [63:0] io_mem0_addr,
  output [63:0] io_mem0_wdata,
  output [7:0]  io_mem0_wmask,
  input         io_mem0_ok,
  input  [63:0] io_mem0_rdata,
  output        io_mem1_en,
  output        io_mem1_op,
  output [63:0] io_mem1_addr,
  output [63:0] io_mem1_wdata,
  output [7:0]  io_mem1_wmask,
  input  [63:0] io_mem1_rdata,
  output        io_mem2_en,
  output        io_mem2_op,
  output [63:0] io_mem2_addr,
  output [63:0] io_mem2_wdata,
  output [7:0]  io_mem2_wmask,
  output [31:0] io_mem2_transfer,
  input         io_mem2_ok,
  input  [63:0] io_mem2_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [1:0] _GEN_0 = io_dmem_addr < 64'h80000000 ? 2'h2 : 2'h0; // @[MMIO.scala 61:48 MMIO.scala 61:53 MMIO.scala 62:24]
  wire [1:0] _GEN_1 = 64'h2000000 <= io_dmem_addr & io_dmem_addr < 64'h200c000 ? 2'h1 : _GEN_0; // @[MMIO.scala 60:76 MMIO.scala 60:81]
  wire [1:0] _GEN_2 = ~io_mem2_ok ? 2'h2 : _GEN_1; // @[MMIO.scala 57:27 MMIO.scala 57:32]
  wire [1:0] sel = ~io_mem0_ok ? 2'h0 : _GEN_2; // @[MMIO.scala 55:22 MMIO.scala 55:27]
  reg [1:0] sel_r; // @[Reg.scala 27:20]
  wire  out_ok = 2'h2 == sel_r ? io_mem2_ok : 2'h1 == sel_r | 2'h0 == sel_r & io_mem0_ok; // @[Mux.scala 80:57]
  wire  _sel_r_T = out_ok & io_dmem_en; // @[MMIO.scala 65:44]
  wire  _io_mem0_en_T = sel == 2'h0; // @[MMIO.scala 67:36]
  wire  _io_mem1_en_T = sel == 2'h1; // @[MMIO.scala 73:36]
  wire  _io_mem2_en_T = sel == 2'h2; // @[MMIO.scala 79:36]
  wire [63:0] _out_rdata_T_1 = 2'h0 == sel_r ? io_mem0_rdata : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _out_rdata_T_3 = 2'h1 == sel_r ? io_mem1_rdata : _out_rdata_T_1; // @[Mux.scala 80:57]
  assign io_dmem_ok = 2'h2 == sel_r ? io_mem2_ok : 2'h1 == sel_r | 2'h0 == sel_r & io_mem0_ok; // @[Mux.scala 80:57]
  assign io_dmem_rdata = 2'h2 == sel_r ? io_mem2_rdata : _out_rdata_T_3; // @[Mux.scala 80:57]
  assign io_mem0_en = sel == 2'h0 & io_dmem_en; // @[MMIO.scala 67:31]
  assign io_mem0_op = _io_mem0_en_T & io_dmem_op; // @[MMIO.scala 68:31]
  assign io_mem0_addr = _io_mem0_en_T ? io_dmem_addr : 64'h0; // @[MMIO.scala 69:31]
  assign io_mem0_wdata = _io_mem0_en_T ? io_dmem_wdata : 64'h0; // @[MMIO.scala 70:31]
  assign io_mem0_wmask = _io_mem0_en_T ? io_dmem_wmask : 8'h0; // @[MMIO.scala 71:31]
  assign io_mem1_en = sel == 2'h1 & io_dmem_en; // @[MMIO.scala 73:31]
  assign io_mem1_op = _io_mem1_en_T & io_dmem_op; // @[MMIO.scala 74:31]
  assign io_mem1_addr = _io_mem1_en_T ? io_dmem_addr : 64'h0; // @[MMIO.scala 75:31]
  assign io_mem1_wdata = _io_mem1_en_T ? io_dmem_wdata : 64'h0; // @[MMIO.scala 76:31]
  assign io_mem1_wmask = _io_mem1_en_T ? io_dmem_wmask : 8'h0; // @[MMIO.scala 77:31]
  assign io_mem2_en = sel == 2'h2 & io_dmem_en; // @[MMIO.scala 79:31]
  assign io_mem2_op = _io_mem2_en_T & io_dmem_op; // @[MMIO.scala 80:31]
  assign io_mem2_addr = _io_mem2_en_T ? io_dmem_addr : 64'h0; // @[MMIO.scala 81:31]
  assign io_mem2_wdata = _io_mem2_en_T ? io_dmem_wdata : 64'h0; // @[MMIO.scala 82:31]
  assign io_mem2_wmask = _io_mem2_en_T ? io_dmem_wmask : 8'h0; // @[MMIO.scala 83:31]
  assign io_mem2_transfer = _io_mem2_en_T ? io_dmem_transfer : 32'h0; // @[MMIO.scala 84:31]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 27:20]
      sel_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_sel_r_T) begin // @[Reg.scala 28:19]
      if (~io_mem0_ok) begin // @[MMIO.scala 55:22]
        sel_r <= 2'h0; // @[MMIO.scala 55:27]
      end else if (~io_mem2_ok) begin // @[MMIO.scala 57:27]
        sel_r <= 2'h2; // @[MMIO.scala 57:32]
      end else begin
        sel_r <= _GEN_1;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sel_r = _RAND_0[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ClintReg(
  input         clock,
  input         reset,
  input         io_mem_en,
  input         io_mem_op,
  input  [63:0] io_mem_addr,
  input  [63:0] io_mem_wdata,
  input  [7:0]  io_mem_wmask,
  output [63:0] io_mem_rdata,
  output        io_set_mtip,
  output        io_clear_mtip
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg  en; // @[MMIO.scala 109:26]
  reg  op; // @[MMIO.scala 110:26]
  reg [63:0] addr; // @[MMIO.scala 111:26]
  reg [63:0] wdata; // @[MMIO.scala 112:26]
  reg [7:0] wm; // @[MMIO.scala 113:26]
  reg [63:0] mtime; // @[MMIO.scala 116:24]
  reg [63:0] mtimecmp; // @[MMIO.scala 117:27]
  wire [7:0] mask64_hi_hi_hi = wm[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] mask64_hi_hi_lo = wm[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] mask64_hi_lo_hi = wm[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] mask64_hi_lo_lo = wm[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] mask64_lo_hi_hi = wm[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] mask64_lo_hi_lo = wm[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] mask64_lo_lo_hi = wm[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] mask64_lo_lo_lo = wm[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [63:0] mask64 = {mask64_hi_hi_hi,mask64_hi_hi_lo,mask64_hi_lo_hi,mask64_hi_lo_lo,mask64_lo_hi_hi,mask64_lo_hi_lo,
    mask64_lo_lo_hi,mask64_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [63:0] _mtime_update_T = ~mask64; // @[MMIO.scala 121:34]
  wire [63:0] _mtime_update_T_1 = mtime & _mtime_update_T; // @[MMIO.scala 121:31]
  wire [63:0] _mtime_update_T_2 = mask64 & wdata; // @[MMIO.scala 121:54]
  wire [63:0] mtime_update = _mtime_update_T_1 | _mtime_update_T_2; // @[MMIO.scala 121:44]
  wire [63:0] _mtimecmp_update_T_1 = mtimecmp & _mtime_update_T; // @[MMIO.scala 122:37]
  wire [63:0] mtimecmp_update = _mtimecmp_update_T_1 | _mtime_update_T_2; // @[MMIO.scala 122:50]
  wire  sel_hi = addr == 64'h2004000; // @[MMIO.scala 124:24]
  wire  sel_lo = addr == 64'h200bff8; // @[MMIO.scala 124:48]
  wire [1:0] sel = {sel_hi,sel_lo}; // @[Cat.scala 30:58]
  wire  _T = en & op; // @[MMIO.scala 134:13]
  wire [63:0] _mtime_T_1 = mtime + 64'h1; // @[MMIO.scala 137:24]
  wire  _T_4 = sel == 2'h2; // @[MMIO.scala 140:26]
  wire [63:0] _io_mem_rdata_T_1 = 2'h1 == sel ? mtime : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _io_mem_rdata_T_3 = 2'h2 == sel ? mtimecmp : _io_mem_rdata_T_1; // @[Mux.scala 80:57]
  assign io_mem_rdata = en & ~op ? _io_mem_rdata_T_3 : 64'h0; // @[MMIO.scala 144:20 MMIO.scala 145:22 MMIO.scala 150:29]
  assign io_set_mtip = ~io_clear_mtip & mtimecmp <= mtime; // @[MMIO.scala 151:35]
  assign io_clear_mtip = _T & _T_4; // @[MMIO.scala 152:31]
  always @(posedge clock) begin
    if (reset) begin // @[MMIO.scala 109:26]
      en <= 1'h0; // @[MMIO.scala 109:26]
    end else begin
      en <= io_mem_en; // @[MMIO.scala 109:26]
    end
    if (reset) begin // @[MMIO.scala 110:26]
      op <= 1'h0; // @[MMIO.scala 110:26]
    end else begin
      op <= io_mem_op; // @[MMIO.scala 110:26]
    end
    if (reset) begin // @[MMIO.scala 111:26]
      addr <= 64'h0; // @[MMIO.scala 111:26]
    end else begin
      addr <= io_mem_addr; // @[MMIO.scala 111:26]
    end
    if (reset) begin // @[MMIO.scala 112:26]
      wdata <= 64'h0; // @[MMIO.scala 112:26]
    end else begin
      wdata <= io_mem_wdata; // @[MMIO.scala 112:26]
    end
    if (reset) begin // @[MMIO.scala 113:26]
      wm <= 8'h0; // @[MMIO.scala 113:26]
    end else begin
      wm <= io_mem_wmask; // @[MMIO.scala 113:26]
    end
    if (reset) begin // @[MMIO.scala 116:24]
      mtime <= 64'h0; // @[MMIO.scala 116:24]
    end else if (en & op & sel == 2'h1) begin // @[MMIO.scala 134:38]
      mtime <= mtime_update; // @[MMIO.scala 134:45]
    end else begin
      mtime <= _mtime_T_1; // @[MMIO.scala 137:15]
    end
    if (reset) begin // @[MMIO.scala 117:27]
      mtimecmp <= 64'h0; // @[MMIO.scala 117:27]
    end else if (_T & sel == 2'h2) begin // @[MMIO.scala 140:38]
      mtimecmp <= mtimecmp_update; // @[MMIO.scala 140:48]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  en = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  op = _RAND_1[0:0];
  _RAND_2 = {2{`RANDOM}};
  addr = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  wdata = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  wm = _RAND_4[7:0];
  _RAND_5 = {2{`RANDOM}};
  mtime = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  mtimecmp = _RAND_6[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DCacheBypass(
  input         clock,
  input         reset,
  input         io_dmem_en,
  input         io_dmem_op,
  input  [63:0] io_dmem_addr,
  input  [63:0] io_dmem_wdata,
  input  [7:0]  io_dmem_wmask,
  input  [31:0] io_dmem_transfer,
  output        io_dmem_ok,
  output [63:0] io_dmem_rdata,
  output        io_axi_req,
  output [31:0] io_axi_raddr,
  input         io_axi_rvalid,
  input  [63:0] io_axi_rdata,
  output        io_axi_weq,
  output [31:0] io_axi_waddr,
  output [63:0] io_axi_wdata,
  output [7:0]  io_axi_wmask,
  input         io_axi_wdone,
  output [2:0]  io_axi_transfer
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] addr; // @[CacheBypass.scala 68:26]
  reg [63:0] wdata; // @[CacheBypass.scala 69:26]
  reg [7:0] wmask; // @[CacheBypass.scala 70:26]
  reg [63:0] rdata; // @[CacheBypass.scala 71:26]
  reg [2:0] transfer; // @[CacheBypass.scala 72:27]
  reg [1:0] state; // @[CacheBypass.scala 75:24]
  wire  _T = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_4 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_5 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_6 = 2'h3 == state; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_3 = io_axi_wdone ? 2'h0 : state; // @[CacheBypass.scala 89:32 CacheBypass.scala 89:39 CacheBypass.scala 75:24]
  wire [1:0] _GEN_4 = _T_6 ? _GEN_3 : state; // @[Conditional.scala 39:67 CacheBypass.scala 75:24]
  wire [63:0] _GEN_9 = state == 2'h0 & io_dmem_en ? io_dmem_addr : {{32'd0}, addr}; // @[CacheBypass.scala 93:39 CacheBypass.scala 95:17 CacheBypass.scala 68:26]
  wire [31:0] _GEN_12 = state == 2'h0 & io_dmem_en ? io_dmem_transfer : {{29'd0}, transfer}; // @[CacheBypass.scala 93:39 CacheBypass.scala 98:18 CacheBypass.scala 72:27]
  wire [38:0] _io_axi_raddr_T = 39'hffffffff << transfer; // @[CacheBypass.scala 103:45]
  wire [38:0] _GEN_13 = {{7'd0}, addr}; // @[CacheBypass.scala 103:29]
  wire [38:0] _io_axi_raddr_T_1 = _GEN_13 & _io_axi_raddr_T; // @[CacheBypass.scala 103:29]
  assign io_dmem_ok = state == 2'h0; // @[CacheBypass.scala 113:30]
  assign io_dmem_rdata = rdata; // @[CacheBypass.scala 112:21]
  assign io_axi_req = state == 2'h1; // @[CacheBypass.scala 102:30]
  assign io_axi_raddr = _io_axi_raddr_T_1[31:0]; // @[CacheBypass.scala 103:21]
  assign io_axi_weq = state == 2'h3; // @[CacheBypass.scala 105:30]
  assign io_axi_waddr = _io_axi_raddr_T_1[31:0]; // @[CacheBypass.scala 106:21]
  assign io_axi_wdata = wdata; // @[CacheBypass.scala 107:21]
  assign io_axi_wmask = wmask; // @[CacheBypass.scala 108:21]
  assign io_axi_transfer = transfer; // @[CacheBypass.scala 110:21]
  always @(posedge clock) begin
    if (reset) begin // @[CacheBypass.scala 68:26]
      addr <= 32'h0; // @[CacheBypass.scala 68:26]
    end else begin
      addr <= _GEN_9[31:0];
    end
    if (reset) begin // @[CacheBypass.scala 69:26]
      wdata <= 64'h0; // @[CacheBypass.scala 69:26]
    end else if (state == 2'h0 & io_dmem_en) begin // @[CacheBypass.scala 93:39]
      wdata <= io_dmem_wdata; // @[CacheBypass.scala 96:17]
    end
    if (reset) begin // @[CacheBypass.scala 70:26]
      wmask <= 8'h0; // @[CacheBypass.scala 70:26]
    end else if (state == 2'h0 & io_dmem_en) begin // @[CacheBypass.scala 93:39]
      wmask <= io_dmem_wmask; // @[CacheBypass.scala 97:17]
    end
    if (reset) begin // @[CacheBypass.scala 71:26]
      rdata <= 64'h0; // @[CacheBypass.scala 71:26]
    end else if (state == 2'h2) begin // @[CacheBypass.scala 100:17]
      rdata <= io_axi_rdata;
    end
    if (reset) begin // @[CacheBypass.scala 72:27]
      transfer <= 3'h0; // @[CacheBypass.scala 72:27]
    end else begin
      transfer <= _GEN_12[2:0];
    end
    if (reset) begin // @[CacheBypass.scala 75:24]
      state <= 2'h0; // @[CacheBypass.scala 75:24]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_dmem_en & ~io_dmem_op) begin // @[CacheBypass.scala 79:45]
        state <= 2'h1; // @[CacheBypass.scala 79:52]
      end else if (io_dmem_en & io_dmem_op) begin // @[CacheBypass.scala 80:49]
        state <= 2'h3; // @[CacheBypass.scala 80:56]
      end
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      if (io_axi_rvalid) begin // @[CacheBypass.scala 83:33]
        state <= 2'h2; // @[CacheBypass.scala 83:40]
      end
    end else if (_T_5) begin // @[Conditional.scala 39:67]
      state <= 2'h0; // @[CacheBypass.scala 86:19]
    end else begin
      state <= _GEN_4;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  addr = _RAND_0[31:0];
  _RAND_1 = {2{`RANDOM}};
  wdata = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  wmask = _RAND_2[7:0];
  _RAND_3 = {2{`RANDOM}};
  rdata = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  transfer = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  state = _RAND_5[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SimTop(
  input         clock,
  input         reset,
  input  [63:0] io_logCtrl_log_begin,
  input  [63:0] io_logCtrl_log_end,
  input  [63:0] io_logCtrl_log_level,
  input         io_perfInfo_clean,
  input         io_perfInfo_dump,
  output        io_uart_out_valid,
  output [7:0]  io_uart_out_ch,
  output        io_uart_in_valid,
  input  [7:0]  io_uart_in_ch,
  input         io_memAXI_0_aw_ready,
  output        io_memAXI_0_aw_valid,
  output [7:0]  io_memAXI_0_aw_bits_len,
  output [2:0]  io_memAXI_0_aw_bits_size,
  output [1:0]  io_memAXI_0_aw_bits_burst,
  output        io_memAXI_0_aw_bits_lock,
  output [3:0]  io_memAXI_0_aw_bits_cache,
  output [3:0]  io_memAXI_0_aw_bits_qos,
  output [63:0] io_memAXI_0_aw_bits_addr,
  output [2:0]  io_memAXI_0_aw_bits_prot,
  output [3:0]  io_memAXI_0_aw_bits_id,
  output [3:0]  io_memAXI_0_aw_bits_user,
  input         io_memAXI_0_w_ready,
  output        io_memAXI_0_w_valid,
  output [63:0] io_memAXI_0_w_bits_data,
  output [7:0]  io_memAXI_0_w_bits_strb,
  output        io_memAXI_0_w_bits_last,
  output        io_memAXI_0_b_ready,
  input         io_memAXI_0_b_valid,
  input  [1:0]  io_memAXI_0_b_bits_resp,
  input  [3:0]  io_memAXI_0_b_bits_id,
  input  [3:0]  io_memAXI_0_b_bits_user,
  input         io_memAXI_0_ar_ready,
  output        io_memAXI_0_ar_valid,
  output [7:0]  io_memAXI_0_ar_bits_len,
  output [2:0]  io_memAXI_0_ar_bits_size,
  output [1:0]  io_memAXI_0_ar_bits_burst,
  output        io_memAXI_0_ar_bits_lock,
  output [3:0]  io_memAXI_0_ar_bits_cache,
  output [3:0]  io_memAXI_0_ar_bits_qos,
  output [63:0] io_memAXI_0_ar_bits_addr,
  output [2:0]  io_memAXI_0_ar_bits_prot,
  output [3:0]  io_memAXI_0_ar_bits_id,
  output [3:0]  io_memAXI_0_ar_bits_user,
  output        io_memAXI_0_r_ready,
  input         io_memAXI_0_r_valid,
  input  [1:0]  io_memAXI_0_r_bits_resp,
  input  [63:0] io_memAXI_0_r_bits_data,
  input         io_memAXI_0_r_bits_last,
  input  [3:0]  io_memAXI_0_r_bits_id,
  input  [3:0]  io_memAXI_0_r_bits_user
);
  wire  core_clock; // @[SimTop.scala 14:20]
  wire  core_reset; // @[SimTop.scala 14:20]
  wire [63:0] core_io_imem_addr; // @[SimTop.scala 14:20]
  wire  core_io_imem_en; // @[SimTop.scala 14:20]
  wire [31:0] core_io_imem_data; // @[SimTop.scala 14:20]
  wire  core_io_imem_ok; // @[SimTop.scala 14:20]
  wire  core_io_dmem_en; // @[SimTop.scala 14:20]
  wire  core_io_dmem_op; // @[SimTop.scala 14:20]
  wire [63:0] core_io_dmem_addr; // @[SimTop.scala 14:20]
  wire [63:0] core_io_dmem_wdata; // @[SimTop.scala 14:20]
  wire [7:0] core_io_dmem_wmask; // @[SimTop.scala 14:20]
  wire [31:0] core_io_dmem_transfer; // @[SimTop.scala 14:20]
  wire  core_io_dmem_ok; // @[SimTop.scala 14:20]
  wire [63:0] core_io_dmem_rdata; // @[SimTop.scala 14:20]
  wire  core_io_set_mtip; // @[SimTop.scala 14:20]
  wire  core_io_clear_mtip; // @[SimTop.scala 14:20]
  wire  core_io_ifence_req; // @[SimTop.scala 14:20]
  wire  core_io_ifence_done; // @[SimTop.scala 14:20]
  wire  core_io_dfence_req; // @[SimTop.scala 14:20]
  wire  core_io_dfence_done; // @[SimTop.scala 14:20]
  wire  icache_clock; // @[SimTop.scala 15:22]
  wire  icache_reset; // @[SimTop.scala 15:22]
  wire [63:0] icache_io_imem_addr; // @[SimTop.scala 15:22]
  wire  icache_io_imem_en; // @[SimTop.scala 15:22]
  wire [31:0] icache_io_imem_data; // @[SimTop.scala 15:22]
  wire  icache_io_imem_ok; // @[SimTop.scala 15:22]
  wire  icache_io_axi_req; // @[SimTop.scala 15:22]
  wire [63:0] icache_io_axi_addr; // @[SimTop.scala 15:22]
  wire  icache_io_axi_valid; // @[SimTop.scala 15:22]
  wire [511:0] icache_io_axi_data; // @[SimTop.scala 15:22]
  wire  icache_io_fence_req; // @[SimTop.scala 15:22]
  wire  icache_io_fence_done; // @[SimTop.scala 15:22]
  wire  dcache_clock; // @[SimTop.scala 16:22]
  wire  dcache_reset; // @[SimTop.scala 16:22]
  wire  dcache_io_dmem_en; // @[SimTop.scala 16:22]
  wire  dcache_io_dmem_op; // @[SimTop.scala 16:22]
  wire [63:0] dcache_io_dmem_addr; // @[SimTop.scala 16:22]
  wire [63:0] dcache_io_dmem_wdata; // @[SimTop.scala 16:22]
  wire [7:0] dcache_io_dmem_wmask; // @[SimTop.scala 16:22]
  wire  dcache_io_dmem_ok; // @[SimTop.scala 16:22]
  wire [63:0] dcache_io_dmem_rdata; // @[SimTop.scala 16:22]
  wire  dcache_io_axi_req; // @[SimTop.scala 16:22]
  wire [63:0] dcache_io_axi_raddr; // @[SimTop.scala 16:22]
  wire  dcache_io_axi_rvalid; // @[SimTop.scala 16:22]
  wire [511:0] dcache_io_axi_rdata; // @[SimTop.scala 16:22]
  wire  dcache_io_axi_weq; // @[SimTop.scala 16:22]
  wire [63:0] dcache_io_axi_waddr; // @[SimTop.scala 16:22]
  wire [511:0] dcache_io_axi_wdata; // @[SimTop.scala 16:22]
  wire  dcache_io_axi_wdone; // @[SimTop.scala 16:22]
  wire  dcache_io_fence_req; // @[SimTop.scala 16:22]
  wire  dcache_io_fence_done; // @[SimTop.scala 16:22]
  wire  axi_clock; // @[SimTop.scala 17:19]
  wire  axi_reset; // @[SimTop.scala 17:19]
  wire  axi_io_out_aw_ready; // @[SimTop.scala 17:19]
  wire  axi_io_out_aw_valid; // @[SimTop.scala 17:19]
  wire [7:0] axi_io_out_aw_bits_len; // @[SimTop.scala 17:19]
  wire [2:0] axi_io_out_aw_bits_size; // @[SimTop.scala 17:19]
  wire [63:0] axi_io_out_aw_bits_addr; // @[SimTop.scala 17:19]
  wire  axi_io_out_w_ready; // @[SimTop.scala 17:19]
  wire  axi_io_out_w_valid; // @[SimTop.scala 17:19]
  wire [63:0] axi_io_out_w_bits_data; // @[SimTop.scala 17:19]
  wire [7:0] axi_io_out_w_bits_strb; // @[SimTop.scala 17:19]
  wire  axi_io_out_w_bits_last; // @[SimTop.scala 17:19]
  wire  axi_io_out_b_ready; // @[SimTop.scala 17:19]
  wire  axi_io_out_b_valid; // @[SimTop.scala 17:19]
  wire  axi_io_out_ar_ready; // @[SimTop.scala 17:19]
  wire  axi_io_out_ar_valid; // @[SimTop.scala 17:19]
  wire [7:0] axi_io_out_ar_bits_len; // @[SimTop.scala 17:19]
  wire [2:0] axi_io_out_ar_bits_size; // @[SimTop.scala 17:19]
  wire [63:0] axi_io_out_ar_bits_addr; // @[SimTop.scala 17:19]
  wire  axi_io_out_r_ready; // @[SimTop.scala 17:19]
  wire  axi_io_out_r_valid; // @[SimTop.scala 17:19]
  wire [63:0] axi_io_out_r_bits_data; // @[SimTop.scala 17:19]
  wire  axi_io_out_r_bits_last; // @[SimTop.scala 17:19]
  wire  axi_io_icacheio_req; // @[SimTop.scala 17:19]
  wire [63:0] axi_io_icacheio_addr; // @[SimTop.scala 17:19]
  wire  axi_io_icacheio_valid; // @[SimTop.scala 17:19]
  wire [511:0] axi_io_icacheio_data; // @[SimTop.scala 17:19]
  wire  axi_io_dcacheio_req; // @[SimTop.scala 17:19]
  wire [63:0] axi_io_dcacheio_raddr; // @[SimTop.scala 17:19]
  wire  axi_io_dcacheio_rvalid; // @[SimTop.scala 17:19]
  wire [511:0] axi_io_dcacheio_rdata; // @[SimTop.scala 17:19]
  wire  axi_io_dcacheio_weq; // @[SimTop.scala 17:19]
  wire [63:0] axi_io_dcacheio_waddr; // @[SimTop.scala 17:19]
  wire [511:0] axi_io_dcacheio_wdata; // @[SimTop.scala 17:19]
  wire  axi_io_dcacheio_wdone; // @[SimTop.scala 17:19]
  wire  axi_io_icacheBypassIO_req; // @[SimTop.scala 17:19]
  wire [31:0] axi_io_icacheBypassIO_addr; // @[SimTop.scala 17:19]
  wire  axi_io_icacheBypassIO_valid; // @[SimTop.scala 17:19]
  wire [63:0] axi_io_icacheBypassIO_data; // @[SimTop.scala 17:19]
  wire  axi_io_dcacheBypassIO_req; // @[SimTop.scala 17:19]
  wire [31:0] axi_io_dcacheBypassIO_raddr; // @[SimTop.scala 17:19]
  wire  axi_io_dcacheBypassIO_rvalid; // @[SimTop.scala 17:19]
  wire [63:0] axi_io_dcacheBypassIO_rdata; // @[SimTop.scala 17:19]
  wire  axi_io_dcacheBypassIO_weq; // @[SimTop.scala 17:19]
  wire [31:0] axi_io_dcacheBypassIO_waddr; // @[SimTop.scala 17:19]
  wire [63:0] axi_io_dcacheBypassIO_wdata; // @[SimTop.scala 17:19]
  wire [7:0] axi_io_dcacheBypassIO_wmask; // @[SimTop.scala 17:19]
  wire  axi_io_dcacheBypassIO_wdone; // @[SimTop.scala 17:19]
  wire [2:0] axi_io_dcacheBypassIO_transfer; // @[SimTop.scala 17:19]
  wire  icacheaxi_clock; // @[SimTop.scala 21:25]
  wire  icacheaxi_reset; // @[SimTop.scala 21:25]
  wire  icacheaxi_io_in_req; // @[SimTop.scala 21:25]
  wire [63:0] icacheaxi_io_in_addr; // @[SimTop.scala 21:25]
  wire  icacheaxi_io_in_valid; // @[SimTop.scala 21:25]
  wire [511:0] icacheaxi_io_in_data; // @[SimTop.scala 21:25]
  wire  icacheaxi_io_out0_req; // @[SimTop.scala 21:25]
  wire [63:0] icacheaxi_io_out0_addr; // @[SimTop.scala 21:25]
  wire  icacheaxi_io_out0_valid; // @[SimTop.scala 21:25]
  wire [511:0] icacheaxi_io_out0_data; // @[SimTop.scala 21:25]
  wire  icacheaxi_io_out1_req; // @[SimTop.scala 21:25]
  wire [31:0] icacheaxi_io_out1_addr; // @[SimTop.scala 21:25]
  wire  icacheaxi_io_out1_valid; // @[SimTop.scala 21:25]
  wire [63:0] icacheaxi_io_out1_data; // @[SimTop.scala 21:25]
  wire  dmmio_clock; // @[SimTop.scala 22:21]
  wire  dmmio_reset; // @[SimTop.scala 22:21]
  wire  dmmio_io_dmem_en; // @[SimTop.scala 22:21]
  wire  dmmio_io_dmem_op; // @[SimTop.scala 22:21]
  wire [63:0] dmmio_io_dmem_addr; // @[SimTop.scala 22:21]
  wire [63:0] dmmio_io_dmem_wdata; // @[SimTop.scala 22:21]
  wire [7:0] dmmio_io_dmem_wmask; // @[SimTop.scala 22:21]
  wire [31:0] dmmio_io_dmem_transfer; // @[SimTop.scala 22:21]
  wire  dmmio_io_dmem_ok; // @[SimTop.scala 22:21]
  wire [63:0] dmmio_io_dmem_rdata; // @[SimTop.scala 22:21]
  wire  dmmio_io_mem0_en; // @[SimTop.scala 22:21]
  wire  dmmio_io_mem0_op; // @[SimTop.scala 22:21]
  wire [63:0] dmmio_io_mem0_addr; // @[SimTop.scala 22:21]
  wire [63:0] dmmio_io_mem0_wdata; // @[SimTop.scala 22:21]
  wire [7:0] dmmio_io_mem0_wmask; // @[SimTop.scala 22:21]
  wire  dmmio_io_mem0_ok; // @[SimTop.scala 22:21]
  wire [63:0] dmmio_io_mem0_rdata; // @[SimTop.scala 22:21]
  wire  dmmio_io_mem1_en; // @[SimTop.scala 22:21]
  wire  dmmio_io_mem1_op; // @[SimTop.scala 22:21]
  wire [63:0] dmmio_io_mem1_addr; // @[SimTop.scala 22:21]
  wire [63:0] dmmio_io_mem1_wdata; // @[SimTop.scala 22:21]
  wire [7:0] dmmio_io_mem1_wmask; // @[SimTop.scala 22:21]
  wire [63:0] dmmio_io_mem1_rdata; // @[SimTop.scala 22:21]
  wire  dmmio_io_mem2_en; // @[SimTop.scala 22:21]
  wire  dmmio_io_mem2_op; // @[SimTop.scala 22:21]
  wire [63:0] dmmio_io_mem2_addr; // @[SimTop.scala 22:21]
  wire [63:0] dmmio_io_mem2_wdata; // @[SimTop.scala 22:21]
  wire [7:0] dmmio_io_mem2_wmask; // @[SimTop.scala 22:21]
  wire [31:0] dmmio_io_mem2_transfer; // @[SimTop.scala 22:21]
  wire  dmmio_io_mem2_ok; // @[SimTop.scala 22:21]
  wire [63:0] dmmio_io_mem2_rdata; // @[SimTop.scala 22:21]
  wire  clintreg_clock; // @[SimTop.scala 23:24]
  wire  clintreg_reset; // @[SimTop.scala 23:24]
  wire  clintreg_io_mem_en; // @[SimTop.scala 23:24]
  wire  clintreg_io_mem_op; // @[SimTop.scala 23:24]
  wire [63:0] clintreg_io_mem_addr; // @[SimTop.scala 23:24]
  wire [63:0] clintreg_io_mem_wdata; // @[SimTop.scala 23:24]
  wire [7:0] clintreg_io_mem_wmask; // @[SimTop.scala 23:24]
  wire [63:0] clintreg_io_mem_rdata; // @[SimTop.scala 23:24]
  wire  clintreg_io_set_mtip; // @[SimTop.scala 23:24]
  wire  clintreg_io_clear_mtip; // @[SimTop.scala 23:24]
  wire  dcachebypass_clock; // @[SimTop.scala 24:28]
  wire  dcachebypass_reset; // @[SimTop.scala 24:28]
  wire  dcachebypass_io_dmem_en; // @[SimTop.scala 24:28]
  wire  dcachebypass_io_dmem_op; // @[SimTop.scala 24:28]
  wire [63:0] dcachebypass_io_dmem_addr; // @[SimTop.scala 24:28]
  wire [63:0] dcachebypass_io_dmem_wdata; // @[SimTop.scala 24:28]
  wire [7:0] dcachebypass_io_dmem_wmask; // @[SimTop.scala 24:28]
  wire [31:0] dcachebypass_io_dmem_transfer; // @[SimTop.scala 24:28]
  wire  dcachebypass_io_dmem_ok; // @[SimTop.scala 24:28]
  wire [63:0] dcachebypass_io_dmem_rdata; // @[SimTop.scala 24:28]
  wire  dcachebypass_io_axi_req; // @[SimTop.scala 24:28]
  wire [31:0] dcachebypass_io_axi_raddr; // @[SimTop.scala 24:28]
  wire  dcachebypass_io_axi_rvalid; // @[SimTop.scala 24:28]
  wire [63:0] dcachebypass_io_axi_rdata; // @[SimTop.scala 24:28]
  wire  dcachebypass_io_axi_weq; // @[SimTop.scala 24:28]
  wire [31:0] dcachebypass_io_axi_waddr; // @[SimTop.scala 24:28]
  wire [63:0] dcachebypass_io_axi_wdata; // @[SimTop.scala 24:28]
  wire [7:0] dcachebypass_io_axi_wmask; // @[SimTop.scala 24:28]
  wire  dcachebypass_io_axi_wdone; // @[SimTop.scala 24:28]
  wire [2:0] dcachebypass_io_axi_transfer; // @[SimTop.scala 24:28]
  Core core ( // @[SimTop.scala 14:20]
    .clock(core_clock),
    .reset(core_reset),
    .io_imem_addr(core_io_imem_addr),
    .io_imem_en(core_io_imem_en),
    .io_imem_data(core_io_imem_data),
    .io_imem_ok(core_io_imem_ok),
    .io_dmem_en(core_io_dmem_en),
    .io_dmem_op(core_io_dmem_op),
    .io_dmem_addr(core_io_dmem_addr),
    .io_dmem_wdata(core_io_dmem_wdata),
    .io_dmem_wmask(core_io_dmem_wmask),
    .io_dmem_transfer(core_io_dmem_transfer),
    .io_dmem_ok(core_io_dmem_ok),
    .io_dmem_rdata(core_io_dmem_rdata),
    .io_set_mtip(core_io_set_mtip),
    .io_clear_mtip(core_io_clear_mtip),
    .io_ifence_req(core_io_ifence_req),
    .io_ifence_done(core_io_ifence_done),
    .io_dfence_req(core_io_dfence_req),
    .io_dfence_done(core_io_dfence_done)
  );
  ICache icache ( // @[SimTop.scala 15:22]
    .clock(icache_clock),
    .reset(icache_reset),
    .io_imem_addr(icache_io_imem_addr),
    .io_imem_en(icache_io_imem_en),
    .io_imem_data(icache_io_imem_data),
    .io_imem_ok(icache_io_imem_ok),
    .io_axi_req(icache_io_axi_req),
    .io_axi_addr(icache_io_axi_addr),
    .io_axi_valid(icache_io_axi_valid),
    .io_axi_data(icache_io_axi_data),
    .io_fence_req(icache_io_fence_req),
    .io_fence_done(icache_io_fence_done)
  );
  DCache dcache ( // @[SimTop.scala 16:22]
    .clock(dcache_clock),
    .reset(dcache_reset),
    .io_dmem_en(dcache_io_dmem_en),
    .io_dmem_op(dcache_io_dmem_op),
    .io_dmem_addr(dcache_io_dmem_addr),
    .io_dmem_wdata(dcache_io_dmem_wdata),
    .io_dmem_wmask(dcache_io_dmem_wmask),
    .io_dmem_ok(dcache_io_dmem_ok),
    .io_dmem_rdata(dcache_io_dmem_rdata),
    .io_axi_req(dcache_io_axi_req),
    .io_axi_raddr(dcache_io_axi_raddr),
    .io_axi_rvalid(dcache_io_axi_rvalid),
    .io_axi_rdata(dcache_io_axi_rdata),
    .io_axi_weq(dcache_io_axi_weq),
    .io_axi_waddr(dcache_io_axi_waddr),
    .io_axi_wdata(dcache_io_axi_wdata),
    .io_axi_wdone(dcache_io_axi_wdone),
    .io_fence_req(dcache_io_fence_req),
    .io_fence_done(dcache_io_fence_done)
  );
  AXI axi ( // @[SimTop.scala 17:19]
    .clock(axi_clock),
    .reset(axi_reset),
    .io_out_aw_ready(axi_io_out_aw_ready),
    .io_out_aw_valid(axi_io_out_aw_valid),
    .io_out_aw_bits_len(axi_io_out_aw_bits_len),
    .io_out_aw_bits_size(axi_io_out_aw_bits_size),
    .io_out_aw_bits_addr(axi_io_out_aw_bits_addr),
    .io_out_w_ready(axi_io_out_w_ready),
    .io_out_w_valid(axi_io_out_w_valid),
    .io_out_w_bits_data(axi_io_out_w_bits_data),
    .io_out_w_bits_strb(axi_io_out_w_bits_strb),
    .io_out_w_bits_last(axi_io_out_w_bits_last),
    .io_out_b_ready(axi_io_out_b_ready),
    .io_out_b_valid(axi_io_out_b_valid),
    .io_out_ar_ready(axi_io_out_ar_ready),
    .io_out_ar_valid(axi_io_out_ar_valid),
    .io_out_ar_bits_len(axi_io_out_ar_bits_len),
    .io_out_ar_bits_size(axi_io_out_ar_bits_size),
    .io_out_ar_bits_addr(axi_io_out_ar_bits_addr),
    .io_out_r_ready(axi_io_out_r_ready),
    .io_out_r_valid(axi_io_out_r_valid),
    .io_out_r_bits_data(axi_io_out_r_bits_data),
    .io_out_r_bits_last(axi_io_out_r_bits_last),
    .io_icacheio_req(axi_io_icacheio_req),
    .io_icacheio_addr(axi_io_icacheio_addr),
    .io_icacheio_valid(axi_io_icacheio_valid),
    .io_icacheio_data(axi_io_icacheio_data),
    .io_dcacheio_req(axi_io_dcacheio_req),
    .io_dcacheio_raddr(axi_io_dcacheio_raddr),
    .io_dcacheio_rvalid(axi_io_dcacheio_rvalid),
    .io_dcacheio_rdata(axi_io_dcacheio_rdata),
    .io_dcacheio_weq(axi_io_dcacheio_weq),
    .io_dcacheio_waddr(axi_io_dcacheio_waddr),
    .io_dcacheio_wdata(axi_io_dcacheio_wdata),
    .io_dcacheio_wdone(axi_io_dcacheio_wdone),
    .io_icacheBypassIO_req(axi_io_icacheBypassIO_req),
    .io_icacheBypassIO_addr(axi_io_icacheBypassIO_addr),
    .io_icacheBypassIO_valid(axi_io_icacheBypassIO_valid),
    .io_icacheBypassIO_data(axi_io_icacheBypassIO_data),
    .io_dcacheBypassIO_req(axi_io_dcacheBypassIO_req),
    .io_dcacheBypassIO_raddr(axi_io_dcacheBypassIO_raddr),
    .io_dcacheBypassIO_rvalid(axi_io_dcacheBypassIO_rvalid),
    .io_dcacheBypassIO_rdata(axi_io_dcacheBypassIO_rdata),
    .io_dcacheBypassIO_weq(axi_io_dcacheBypassIO_weq),
    .io_dcacheBypassIO_waddr(axi_io_dcacheBypassIO_waddr),
    .io_dcacheBypassIO_wdata(axi_io_dcacheBypassIO_wdata),
    .io_dcacheBypassIO_wmask(axi_io_dcacheBypassIO_wmask),
    .io_dcacheBypassIO_wdone(axi_io_dcacheBypassIO_wdone),
    .io_dcacheBypassIO_transfer(axi_io_dcacheBypassIO_transfer)
  );
  ICacheSocAxi icacheaxi ( // @[SimTop.scala 21:25]
    .clock(icacheaxi_clock),
    .reset(icacheaxi_reset),
    .io_in_req(icacheaxi_io_in_req),
    .io_in_addr(icacheaxi_io_in_addr),
    .io_in_valid(icacheaxi_io_in_valid),
    .io_in_data(icacheaxi_io_in_data),
    .io_out0_req(icacheaxi_io_out0_req),
    .io_out0_addr(icacheaxi_io_out0_addr),
    .io_out0_valid(icacheaxi_io_out0_valid),
    .io_out0_data(icacheaxi_io_out0_data),
    .io_out1_req(icacheaxi_io_out1_req),
    .io_out1_addr(icacheaxi_io_out1_addr),
    .io_out1_valid(icacheaxi_io_out1_valid),
    .io_out1_data(icacheaxi_io_out1_data)
  );
  DMMIO dmmio ( // @[SimTop.scala 22:21]
    .clock(dmmio_clock),
    .reset(dmmio_reset),
    .io_dmem_en(dmmio_io_dmem_en),
    .io_dmem_op(dmmio_io_dmem_op),
    .io_dmem_addr(dmmio_io_dmem_addr),
    .io_dmem_wdata(dmmio_io_dmem_wdata),
    .io_dmem_wmask(dmmio_io_dmem_wmask),
    .io_dmem_transfer(dmmio_io_dmem_transfer),
    .io_dmem_ok(dmmio_io_dmem_ok),
    .io_dmem_rdata(dmmio_io_dmem_rdata),
    .io_mem0_en(dmmio_io_mem0_en),
    .io_mem0_op(dmmio_io_mem0_op),
    .io_mem0_addr(dmmio_io_mem0_addr),
    .io_mem0_wdata(dmmio_io_mem0_wdata),
    .io_mem0_wmask(dmmio_io_mem0_wmask),
    .io_mem0_ok(dmmio_io_mem0_ok),
    .io_mem0_rdata(dmmio_io_mem0_rdata),
    .io_mem1_en(dmmio_io_mem1_en),
    .io_mem1_op(dmmio_io_mem1_op),
    .io_mem1_addr(dmmio_io_mem1_addr),
    .io_mem1_wdata(dmmio_io_mem1_wdata),
    .io_mem1_wmask(dmmio_io_mem1_wmask),
    .io_mem1_rdata(dmmio_io_mem1_rdata),
    .io_mem2_en(dmmio_io_mem2_en),
    .io_mem2_op(dmmio_io_mem2_op),
    .io_mem2_addr(dmmio_io_mem2_addr),
    .io_mem2_wdata(dmmio_io_mem2_wdata),
    .io_mem2_wmask(dmmio_io_mem2_wmask),
    .io_mem2_transfer(dmmio_io_mem2_transfer),
    .io_mem2_ok(dmmio_io_mem2_ok),
    .io_mem2_rdata(dmmio_io_mem2_rdata)
  );
  ClintReg clintreg ( // @[SimTop.scala 23:24]
    .clock(clintreg_clock),
    .reset(clintreg_reset),
    .io_mem_en(clintreg_io_mem_en),
    .io_mem_op(clintreg_io_mem_op),
    .io_mem_addr(clintreg_io_mem_addr),
    .io_mem_wdata(clintreg_io_mem_wdata),
    .io_mem_wmask(clintreg_io_mem_wmask),
    .io_mem_rdata(clintreg_io_mem_rdata),
    .io_set_mtip(clintreg_io_set_mtip),
    .io_clear_mtip(clintreg_io_clear_mtip)
  );
  DCacheBypass dcachebypass ( // @[SimTop.scala 24:28]
    .clock(dcachebypass_clock),
    .reset(dcachebypass_reset),
    .io_dmem_en(dcachebypass_io_dmem_en),
    .io_dmem_op(dcachebypass_io_dmem_op),
    .io_dmem_addr(dcachebypass_io_dmem_addr),
    .io_dmem_wdata(dcachebypass_io_dmem_wdata),
    .io_dmem_wmask(dcachebypass_io_dmem_wmask),
    .io_dmem_transfer(dcachebypass_io_dmem_transfer),
    .io_dmem_ok(dcachebypass_io_dmem_ok),
    .io_dmem_rdata(dcachebypass_io_dmem_rdata),
    .io_axi_req(dcachebypass_io_axi_req),
    .io_axi_raddr(dcachebypass_io_axi_raddr),
    .io_axi_rvalid(dcachebypass_io_axi_rvalid),
    .io_axi_rdata(dcachebypass_io_axi_rdata),
    .io_axi_weq(dcachebypass_io_axi_weq),
    .io_axi_waddr(dcachebypass_io_axi_waddr),
    .io_axi_wdata(dcachebypass_io_axi_wdata),
    .io_axi_wmask(dcachebypass_io_axi_wmask),
    .io_axi_wdone(dcachebypass_io_axi_wdone),
    .io_axi_transfer(dcachebypass_io_axi_transfer)
  );
  assign io_uart_out_valid = 1'h0; // @[SimTop.scala 52:21]
  assign io_uart_out_ch = 8'h0; // @[SimTop.scala 53:18]
  assign io_uart_in_valid = 1'h0; // @[SimTop.scala 54:20]
  assign io_memAXI_0_aw_valid = axi_io_out_aw_valid; // @[SimTop.scala 48:17]
  assign io_memAXI_0_aw_bits_len = axi_io_out_aw_bits_len; // @[SimTop.scala 48:17]
  assign io_memAXI_0_aw_bits_size = axi_io_out_aw_bits_size; // @[SimTop.scala 48:17]
  assign io_memAXI_0_aw_bits_burst = 2'h1; // @[SimTop.scala 48:17]
  assign io_memAXI_0_aw_bits_lock = 1'h0; // @[SimTop.scala 48:17]
  assign io_memAXI_0_aw_bits_cache = 4'h2; // @[SimTop.scala 48:17]
  assign io_memAXI_0_aw_bits_qos = 4'h0; // @[SimTop.scala 48:17]
  assign io_memAXI_0_aw_bits_addr = axi_io_out_aw_bits_addr; // @[SimTop.scala 48:17]
  assign io_memAXI_0_aw_bits_prot = 3'h0; // @[SimTop.scala 48:17]
  assign io_memAXI_0_aw_bits_id = 4'h0; // @[SimTop.scala 48:17]
  assign io_memAXI_0_aw_bits_user = 4'h0; // @[SimTop.scala 48:17]
  assign io_memAXI_0_w_valid = axi_io_out_w_valid; // @[SimTop.scala 49:17]
  assign io_memAXI_0_w_bits_data = axi_io_out_w_bits_data; // @[SimTop.scala 49:17]
  assign io_memAXI_0_w_bits_strb = axi_io_out_w_bits_strb; // @[SimTop.scala 49:17]
  assign io_memAXI_0_w_bits_last = axi_io_out_w_bits_last; // @[SimTop.scala 49:17]
  assign io_memAXI_0_b_ready = axi_io_out_b_ready; // @[SimTop.scala 50:17]
  assign io_memAXI_0_ar_valid = axi_io_out_ar_valid; // @[SimTop.scala 46:17]
  assign io_memAXI_0_ar_bits_len = axi_io_out_ar_bits_len; // @[SimTop.scala 46:17]
  assign io_memAXI_0_ar_bits_size = axi_io_out_ar_bits_size; // @[SimTop.scala 46:17]
  assign io_memAXI_0_ar_bits_burst = 2'h1; // @[SimTop.scala 46:17]
  assign io_memAXI_0_ar_bits_lock = 1'h0; // @[SimTop.scala 46:17]
  assign io_memAXI_0_ar_bits_cache = 4'h2; // @[SimTop.scala 46:17]
  assign io_memAXI_0_ar_bits_qos = 4'h0; // @[SimTop.scala 46:17]
  assign io_memAXI_0_ar_bits_addr = axi_io_out_ar_bits_addr; // @[SimTop.scala 46:17]
  assign io_memAXI_0_ar_bits_prot = 3'h0; // @[SimTop.scala 46:17]
  assign io_memAXI_0_ar_bits_id = 4'h0; // @[SimTop.scala 46:17]
  assign io_memAXI_0_ar_bits_user = 4'h0; // @[SimTop.scala 46:17]
  assign io_memAXI_0_r_ready = axi_io_out_r_ready; // @[SimTop.scala 47:17]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_imem_data = icache_io_imem_data; // @[SimTop.scala 29:17]
  assign core_io_imem_ok = icache_io_imem_ok; // @[SimTop.scala 29:17]
  assign core_io_dmem_ok = dmmio_io_dmem_ok; // @[SimTop.scala 31:17]
  assign core_io_dmem_rdata = dmmio_io_dmem_rdata; // @[SimTop.scala 31:17]
  assign core_io_set_mtip = clintreg_io_set_mtip; // @[SimTop.scala 36:23]
  assign core_io_clear_mtip = clintreg_io_clear_mtip; // @[SimTop.scala 37:23]
  assign core_io_ifence_done = icache_io_fence_done; // @[SimTop.scala 26:19]
  assign core_io_dfence_done = dcache_io_fence_done; // @[SimTop.scala 27:19]
  assign icache_clock = clock;
  assign icache_reset = reset;
  assign icache_io_imem_addr = core_io_imem_addr; // @[SimTop.scala 29:17]
  assign icache_io_imem_en = core_io_imem_en; // @[SimTop.scala 29:17]
  assign icache_io_axi_valid = icacheaxi_io_in_valid; // @[SimTop.scala 39:17]
  assign icache_io_axi_data = icacheaxi_io_in_data; // @[SimTop.scala 39:17]
  assign icache_io_fence_req = core_io_ifence_req; // @[SimTop.scala 26:19]
  assign dcache_clock = clock;
  assign dcache_reset = reset;
  assign dcache_io_dmem_en = dmmio_io_mem0_en; // @[SimTop.scala 32:17]
  assign dcache_io_dmem_op = dmmio_io_mem0_op; // @[SimTop.scala 32:17]
  assign dcache_io_dmem_addr = dmmio_io_mem0_addr; // @[SimTop.scala 32:17]
  assign dcache_io_dmem_wdata = dmmio_io_mem0_wdata; // @[SimTop.scala 32:17]
  assign dcache_io_dmem_wmask = dmmio_io_mem0_wmask; // @[SimTop.scala 32:17]
  assign dcache_io_axi_rvalid = axi_io_dcacheio_rvalid; // @[SimTop.scala 43:17]
  assign dcache_io_axi_rdata = axi_io_dcacheio_rdata; // @[SimTop.scala 43:17]
  assign dcache_io_axi_wdone = axi_io_dcacheio_wdone; // @[SimTop.scala 43:17]
  assign dcache_io_fence_req = core_io_dfence_req; // @[SimTop.scala 27:19]
  assign axi_clock = clock;
  assign axi_reset = reset;
  assign axi_io_out_aw_ready = io_memAXI_0_aw_ready; // @[SimTop.scala 48:17]
  assign axi_io_out_w_ready = io_memAXI_0_w_ready; // @[SimTop.scala 49:17]
  assign axi_io_out_b_valid = io_memAXI_0_b_valid; // @[SimTop.scala 50:17]
  assign axi_io_out_ar_ready = io_memAXI_0_ar_ready; // @[SimTop.scala 46:17]
  assign axi_io_out_r_valid = io_memAXI_0_r_valid; // @[SimTop.scala 47:17]
  assign axi_io_out_r_bits_data = io_memAXI_0_r_bits_data; // @[SimTop.scala 47:17]
  assign axi_io_out_r_bits_last = io_memAXI_0_r_bits_last; // @[SimTop.scala 47:17]
  assign axi_io_icacheio_req = icacheaxi_io_out0_req; // @[SimTop.scala 40:21]
  assign axi_io_icacheio_addr = icacheaxi_io_out0_addr; // @[SimTop.scala 40:21]
  assign axi_io_dcacheio_req = dcache_io_axi_req; // @[SimTop.scala 43:17]
  assign axi_io_dcacheio_raddr = dcache_io_axi_raddr; // @[SimTop.scala 43:17]
  assign axi_io_dcacheio_weq = dcache_io_axi_weq; // @[SimTop.scala 43:17]
  assign axi_io_dcacheio_waddr = dcache_io_axi_waddr; // @[SimTop.scala 43:17]
  assign axi_io_dcacheio_wdata = dcache_io_axi_wdata; // @[SimTop.scala 43:17]
  assign axi_io_icacheBypassIO_req = icacheaxi_io_out1_req; // @[SimTop.scala 41:21]
  assign axi_io_icacheBypassIO_addr = icacheaxi_io_out1_addr; // @[SimTop.scala 41:21]
  assign axi_io_dcacheBypassIO_req = dcachebypass_io_axi_req; // @[SimTop.scala 44:23]
  assign axi_io_dcacheBypassIO_raddr = dcachebypass_io_axi_raddr; // @[SimTop.scala 44:23]
  assign axi_io_dcacheBypassIO_weq = dcachebypass_io_axi_weq; // @[SimTop.scala 44:23]
  assign axi_io_dcacheBypassIO_waddr = dcachebypass_io_axi_waddr; // @[SimTop.scala 44:23]
  assign axi_io_dcacheBypassIO_wdata = dcachebypass_io_axi_wdata; // @[SimTop.scala 44:23]
  assign axi_io_dcacheBypassIO_wmask = dcachebypass_io_axi_wmask; // @[SimTop.scala 44:23]
  assign axi_io_dcacheBypassIO_transfer = dcachebypass_io_axi_transfer; // @[SimTop.scala 44:23]
  assign icacheaxi_clock = clock;
  assign icacheaxi_reset = reset;
  assign icacheaxi_io_in_req = icache_io_axi_req; // @[SimTop.scala 39:17]
  assign icacheaxi_io_in_addr = icache_io_axi_addr; // @[SimTop.scala 39:17]
  assign icacheaxi_io_out0_valid = axi_io_icacheio_valid; // @[SimTop.scala 40:21]
  assign icacheaxi_io_out0_data = axi_io_icacheio_data; // @[SimTop.scala 40:21]
  assign icacheaxi_io_out1_valid = axi_io_icacheBypassIO_valid; // @[SimTop.scala 41:21]
  assign icacheaxi_io_out1_data = axi_io_icacheBypassIO_data; // @[SimTop.scala 41:21]
  assign dmmio_clock = clock;
  assign dmmio_reset = reset;
  assign dmmio_io_dmem_en = core_io_dmem_en; // @[SimTop.scala 31:17]
  assign dmmio_io_dmem_op = core_io_dmem_op; // @[SimTop.scala 31:17]
  assign dmmio_io_dmem_addr = core_io_dmem_addr; // @[SimTop.scala 31:17]
  assign dmmio_io_dmem_wdata = core_io_dmem_wdata; // @[SimTop.scala 31:17]
  assign dmmio_io_dmem_wmask = core_io_dmem_wmask; // @[SimTop.scala 31:17]
  assign dmmio_io_dmem_transfer = core_io_dmem_transfer; // @[SimTop.scala 31:17]
  assign dmmio_io_mem0_ok = dcache_io_dmem_ok; // @[SimTop.scala 32:17]
  assign dmmio_io_mem0_rdata = dcache_io_dmem_rdata; // @[SimTop.scala 32:17]
  assign dmmio_io_mem1_rdata = clintreg_io_mem_rdata; // @[SimTop.scala 33:17]
  assign dmmio_io_mem2_ok = dcachebypass_io_dmem_ok; // @[SimTop.scala 34:17]
  assign dmmio_io_mem2_rdata = dcachebypass_io_dmem_rdata; // @[SimTop.scala 34:17]
  assign clintreg_clock = clock;
  assign clintreg_reset = reset;
  assign clintreg_io_mem_en = dmmio_io_mem1_en; // @[SimTop.scala 33:17]
  assign clintreg_io_mem_op = dmmio_io_mem1_op; // @[SimTop.scala 33:17]
  assign clintreg_io_mem_addr = dmmio_io_mem1_addr; // @[SimTop.scala 33:17]
  assign clintreg_io_mem_wdata = dmmio_io_mem1_wdata; // @[SimTop.scala 33:17]
  assign clintreg_io_mem_wmask = dmmio_io_mem1_wmask; // @[SimTop.scala 33:17]
  assign dcachebypass_clock = clock;
  assign dcachebypass_reset = reset;
  assign dcachebypass_io_dmem_en = dmmio_io_mem2_en; // @[SimTop.scala 34:17]
  assign dcachebypass_io_dmem_op = dmmio_io_mem2_op; // @[SimTop.scala 34:17]
  assign dcachebypass_io_dmem_addr = dmmio_io_mem2_addr; // @[SimTop.scala 34:17]
  assign dcachebypass_io_dmem_wdata = dmmio_io_mem2_wdata; // @[SimTop.scala 34:17]
  assign dcachebypass_io_dmem_wmask = dmmio_io_mem2_wmask; // @[SimTop.scala 34:17]
  assign dcachebypass_io_dmem_transfer = dmmio_io_mem2_transfer; // @[SimTop.scala 34:17]
  assign dcachebypass_io_axi_rvalid = axi_io_dcacheBypassIO_rvalid; // @[SimTop.scala 44:23]
  assign dcachebypass_io_axi_rdata = axi_io_dcacheBypassIO_rdata; // @[SimTop.scala 44:23]
  assign dcachebypass_io_axi_wdone = axi_io_dcacheBypassIO_wdone; // @[SimTop.scala 44:23]
endmodule
