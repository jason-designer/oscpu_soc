module IFetch(
  input         reset,
  input         io_jump_en,
  input  [63:0] io_jump_pc,
  input         io_en,
  input  [63:0] io_pc,
  output [63:0] io_next_pc,
  output        io_valid
);
  wire [63:0] _io_next_pc_T_1 = io_pc + 64'h4; // @[IFetch.scala 14:69]
  wire [63:0] _io_next_pc_T_2 = io_jump_en ? io_jump_pc : _io_next_pc_T_1; // @[IFetch.scala 14:38]
  assign io_next_pc = io_en ? io_pc : _io_next_pc_T_2; // @[IFetch.scala 14:20]
  assign io_valid = ~reset; // @[IFetch.scala 15:17]
endmodule
module Decode(
  input  [63:0] io_pc,
  input  [31:0] io_inst,
  output        io_rs1_en,
  output        io_rs2_en,
  output [4:0]  io_rs1_addr,
  output [4:0]  io_rs2_addr,
  input  [63:0] io_rs1_data,
  input  [63:0] io_rs2_data,
  output        io_rd_en,
  output [4:0]  io_rd_addr,
  output [5:0]  io_decode_info_fu_code,
  output [15:0] io_decode_info_alu_code,
  output [7:0]  io_decode_info_bu_code,
  output [6:0]  io_decode_info_lu_code,
  output [3:0]  io_decode_info_su_code,
  output [9:0]  io_decode_info_mdu_code,
  output [6:0]  io_decode_info_csru_code,
  output        io_jump_en,
  output [63:0] io_jump_pc,
  output [63:0] io_op1,
  output [63:0] io_op2,
  output [63:0] io_imm,
  output        io_putch,
  input  [63:0] io_mtvec,
  input  [63:0] io_mepc
);
  wire [31:0] _sll_T = io_inst & 32'hfe00707f; // @[Decode.scala 47:20]
  wire  sll = 32'h1033 == _sll_T; // @[Decode.scala 47:20]
  wire  srl = 32'h5033 == _sll_T; // @[Decode.scala 48:20]
  wire  sra = 32'h40005033 == _sll_T; // @[Decode.scala 49:20]
  wire [31:0] _slli_T = io_inst & 32'hfc00707f; // @[Decode.scala 50:21]
  wire  slli = 32'h1013 == _slli_T; // @[Decode.scala 50:21]
  wire  srli = 32'h5013 == _slli_T; // @[Decode.scala 51:21]
  wire  srai = 32'h40005013 == _slli_T; // @[Decode.scala 52:21]
  wire  sllw = 32'h103b == _sll_T; // @[Decode.scala 53:21]
  wire  srlw = 32'h503b == _sll_T; // @[Decode.scala 54:21]
  wire  sraw = 32'h4000503b == _sll_T; // @[Decode.scala 55:21]
  wire  slliw = 32'h101b == _sll_T; // @[Decode.scala 56:22]
  wire  srliw = 32'h501b == _sll_T; // @[Decode.scala 57:22]
  wire  sraiw = 32'h4000501b == _sll_T; // @[Decode.scala 58:22]
  wire  add = 32'h33 == _sll_T; // @[Decode.scala 60:24]
  wire  addw = 32'h3b == _sll_T; // @[Decode.scala 61:24]
  wire [31:0] _addi_T = io_inst & 32'h707f; // @[Decode.scala 62:24]
  wire  addi = 32'h13 == _addi_T; // @[Decode.scala 62:24]
  wire  addiw = 32'h1b == _addi_T; // @[Decode.scala 63:24]
  wire  alu_sub = 32'h40000033 == _sll_T; // @[Decode.scala 64:24]
  wire  alu_subw = 32'h4000003b == _sll_T; // @[Decode.scala 65:24]
  wire [31:0] _lui_T = io_inst & 32'h7f; // @[Decode.scala 66:24]
  wire  lui = 32'h37 == _lui_T; // @[Decode.scala 66:24]
  wire  alu_auipc = 32'h17 == _lui_T; // @[Decode.scala 67:24]
  wire  xor_ = 32'h4033 == _sll_T; // @[Decode.scala 69:24]
  wire  or_ = 32'h6033 == _sll_T; // @[Decode.scala 70:24]
  wire  and_ = 32'h7033 == _sll_T; // @[Decode.scala 71:24]
  wire  xori = 32'h4013 == _addi_T; // @[Decode.scala 72:24]
  wire  ori = 32'h6013 == _addi_T; // @[Decode.scala 73:24]
  wire  andi = 32'h7013 == _addi_T; // @[Decode.scala 74:24]
  wire  slt = 32'h2033 == _sll_T; // @[Decode.scala 76:24]
  wire  sltu = 32'h3033 == _sll_T; // @[Decode.scala 77:24]
  wire  slti = 32'h2013 == _addi_T; // @[Decode.scala 78:24]
  wire  sltiu = 32'h3013 == _addi_T; // @[Decode.scala 79:24]
  wire  beq = 32'h63 == _addi_T; // @[Decode.scala 81:24]
  wire  bne = 32'h1063 == _addi_T; // @[Decode.scala 82:24]
  wire  blt = 32'h4063 == _addi_T; // @[Decode.scala 83:24]
  wire  bge = 32'h5063 == _addi_T; // @[Decode.scala 84:24]
  wire  bltu = 32'h6063 == _addi_T; // @[Decode.scala 85:24]
  wire  bgeu = 32'h7063 == _addi_T; // @[Decode.scala 86:24]
  wire  jal = 32'h6f == _lui_T; // @[Decode.scala 88:24]
  wire  jalr = 32'h67 == _addi_T; // @[Decode.scala 89:24]
  wire  lb = 32'h3 == _addi_T; // @[Decode.scala 91:24]
  wire  lh = 32'h1003 == _addi_T; // @[Decode.scala 92:24]
  wire  lw = 32'h2003 == _addi_T; // @[Decode.scala 93:24]
  wire  ld = 32'h3003 == _addi_T; // @[Decode.scala 94:24]
  wire  lbu = 32'h4003 == _addi_T; // @[Decode.scala 95:24]
  wire  lhu = 32'h5003 == _addi_T; // @[Decode.scala 96:24]
  wire  lwu = 32'h6003 == _addi_T; // @[Decode.scala 97:24]
  wire  sb = 32'h23 == _addi_T; // @[Decode.scala 99:24]
  wire  sh = 32'h1023 == _addi_T; // @[Decode.scala 100:24]
  wire  sw = 32'h2023 == _addi_T; // @[Decode.scala 101:24]
  wire  sd = 32'h3023 == _addi_T; // @[Decode.scala 102:24]
  wire  mul = 32'h2000033 == _sll_T; // @[Decode.scala 104:24]
  wire  mulw = 32'h200003b == _sll_T; // @[Decode.scala 105:24]
  wire  div = 32'h2004033 == _sll_T; // @[Decode.scala 106:24]
  wire  divw = 32'h200403b == _sll_T; // @[Decode.scala 107:24]
  wire  divu = 32'h2005033 == _sll_T; // @[Decode.scala 108:24]
  wire  divuw = 32'h200503b == _sll_T; // @[Decode.scala 109:24]
  wire  rem = 32'h2006033 == _sll_T; // @[Decode.scala 110:24]
  wire  remw = 32'h200603b == _sll_T; // @[Decode.scala 111:24]
  wire  remu = 32'h2007033 == _sll_T; // @[Decode.scala 112:24]
  wire  remuw = 32'h200703b == _sll_T; // @[Decode.scala 113:24]
  wire  ecall = 32'h73 == io_inst; // @[Decode.scala 115:24]
  wire  mret = 32'h30200073 == io_inst; // @[Decode.scala 116:24]
  wire  csrrs = 32'h2073 == _addi_T; // @[Decode.scala 117:24]
  wire  csrrw = 32'h1073 == _addi_T; // @[Decode.scala 118:24]
  wire  csrrc = 32'h3073 == _addi_T; // @[Decode.scala 119:24]
  wire  csrrwi = 32'h5073 == _addi_T; // @[Decode.scala 120:24]
  wire  csrrci = 32'h7073 == _addi_T; // @[Decode.scala 121:24]
  wire  alu_add = add | addi | lui; // @[Decode.scala 129:33]
  wire  alu_addw = addw | addiw; // @[Decode.scala 130:26]
  wire  alu_sll = sll | slli; // @[Decode.scala 135:26]
  wire  alu_srl = srl | srli; // @[Decode.scala 136:26]
  wire  alu_sra = sra | srai; // @[Decode.scala 137:26]
  wire  alu_sllw = sllw | slliw; // @[Decode.scala 138:26]
  wire  alu_srlw = srlw | srliw; // @[Decode.scala 139:26]
  wire  alu_sraw = sraw | sraiw; // @[Decode.scala 140:26]
  wire  alu_xor = xor_ | xori; // @[Decode.scala 142:26]
  wire  alu_or = or_ | ori; // @[Decode.scala 143:26]
  wire  alu_and = and_ | andi; // @[Decode.scala 144:26]
  wire  alu_slt = slt | slti; // @[Decode.scala 146:26]
  wire  alu_sltu = sltu | sltiu; // @[Decode.scala 147:26]
  wire [7:0] alu_code_lo = {alu_sra,alu_srl,alu_sll,alu_auipc,alu_subw,alu_sub,alu_addw,alu_add}; // @[Cat.scala 30:58]
  wire [7:0] alu_code_hi = {alu_sltu,alu_slt,alu_and,alu_or,alu_xor,alu_sraw,alu_srlw,alu_sllw}; // @[Cat.scala 30:58]
  wire [15:0] alu_code = {alu_sltu,alu_slt,alu_and,alu_or,alu_xor,alu_sraw,alu_srlw,alu_sllw,alu_code_lo}; // @[Cat.scala 30:58]
  wire  alu_en = alu_code != 16'h0; // @[Decode.scala 150:29]
  wire [3:0] bu_code_lo = {bge,blt,bne,beq}; // @[Cat.scala 30:58]
  wire [3:0] bu_code_hi = {jalr,jal,bgeu,bltu}; // @[Cat.scala 30:58]
  wire [7:0] bu_code = {jalr,jal,bgeu,bltu,bge,blt,bne,beq}; // @[Cat.scala 30:58]
  wire  bu_en = bu_code != 8'h0; // @[Decode.scala 153:27]
  wire [2:0] lu_code_lo = {lw,lh,lb}; // @[Cat.scala 30:58]
  wire [3:0] lu_code_hi = {lwu,lhu,lbu,ld}; // @[Cat.scala 30:58]
  wire [6:0] lu_code = {lwu,lhu,lbu,ld,lw,lh,lb}; // @[Cat.scala 30:58]
  wire  lu_en = lu_code != 7'h0; // @[Decode.scala 156:27]
  wire [1:0] su_code_lo = {sh,sb}; // @[Cat.scala 30:58]
  wire [1:0] su_code_hi = {sd,sw}; // @[Cat.scala 30:58]
  wire [3:0] su_code = {sd,sw,sh,sb}; // @[Cat.scala 30:58]
  wire  su_en = su_code != 4'h0; // @[Decode.scala 159:27]
  wire [4:0] mdu_code_lo = {divu,divw,div,mulw,mul}; // @[Cat.scala 30:58]
  wire [4:0] mdu_code_hi = {remuw,remu,remw,rem,divuw}; // @[Cat.scala 30:58]
  wire [9:0] mdu_code = {remuw,remu,remw,rem,divuw,divu,divw,div,mulw,mul}; // @[Cat.scala 30:58]
  wire  mdu_en = mdu_code != 10'h0; // @[Decode.scala 162:29]
  wire [2:0] csru_code_lo = {csrrs,mret,ecall}; // @[Cat.scala 30:58]
  wire [3:0] csru_code_hi = {csrrci,csrrwi,csrrc,csrrw}; // @[Cat.scala 30:58]
  wire [6:0] csru_code = {csrrci,csrrwi,csrrc,csrrw,csrrs,mret,ecall}; // @[Cat.scala 30:58]
  wire  csr_en = csru_code != 7'h0; // @[Decode.scala 165:31]
  wire [2:0] fu_code_lo = {lu_en,bu_en,alu_en}; // @[Cat.scala 30:58]
  wire [2:0] fu_code_hi = {csr_en,mdu_en,su_en}; // @[Cat.scala 30:58]
  wire  _type_r_T_5 = sll | srl | sra | sllw | srlw | sraw | add; // @[Decode.scala 170:74]
  wire  _type_r_T_9 = _type_r_T_5 | addw | alu_sub | alu_subw | xor_; // @[Decode.scala 171:54]
  wire  _type_r_T_12 = _type_r_T_9 | or_ | and_ | slt; // @[Decode.scala 172:45]
  wire  _type_r_T_14 = _type_r_T_12 | sltu | mul; // @[Decode.scala 173:36]
  wire  _type_r_T_16 = _type_r_T_14 | mulw | div; // @[Decode.scala 174:36]
  wire  _type_r_T_20 = _type_r_T_16 | divw | divu | divuw | rem; // @[Decode.scala 175:54]
  wire  type_r = _type_r_T_20 | remw | remu | remuw | mret; // @[Decode.scala 176:54]
  wire  _type_i_T_5 = slli | srli | srai | slliw | srliw | sraiw | addi; // @[Decode.scala 178:74]
  wire  _type_i_T_7 = _type_i_T_5 | addiw | xori; // @[Decode.scala 179:36]
  wire  _type_i_T_10 = _type_i_T_7 | ori | andi | slti; // @[Decode.scala 180:45]
  wire  _type_i_T_12 = _type_i_T_10 | sltiu | jalr; // @[Decode.scala 181:36]
  wire  _type_i_T_13 = _type_i_T_12 | lb; // @[Decode.scala 182:27]
  wire  _type_i_T_20 = _type_i_T_13 | lh | lw | ld | lbu | lhu | lwu | ecall; // @[Decode.scala 183:81]
  wire  type_i = _type_i_T_20 | csrrs | csrrw | csrrc | csrrwi | csrrci; // @[Decode.scala 184:64]
  wire  type_s = sb | sh | sw | sd; // @[Decode.scala 185:45]
  wire  type_b = beq | bne | blt | bge | bltu | bgeu; // @[Decode.scala 186:64]
  wire  type_u = lui | alu_auipc; // @[Decode.scala 187:27]
  wire [5:0] inst_type = {type_r,type_i,type_s,type_b,type_u,jal}; // @[Cat.scala 30:58]
  wire [51:0] imm_i_hi = io_inst[31] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 72:12]
  wire [11:0] imm_i_lo = io_inst[31:20]; // @[Decode.scala 193:45]
  wire [63:0] imm_i = {imm_i_hi,imm_i_lo}; // @[Cat.scala 30:58]
  wire [6:0] imm_s_hi_lo = io_inst[31:25]; // @[Decode.scala 194:45]
  wire [4:0] imm_s_lo = io_inst[11:7]; // @[Decode.scala 194:59]
  wire [63:0] imm_s = {imm_i_hi,imm_s_hi_lo,imm_s_lo}; // @[Cat.scala 30:58]
  wire [50:0] imm_b_hi_hi_hi = io_inst[31] ? 51'h7ffffffffffff : 51'h0; // @[Bitwise.scala 72:12]
  wire  imm_b_hi_lo = io_inst[7]; // @[Decode.scala 195:55]
  wire [5:0] imm_b_lo_hi_hi = io_inst[30:25]; // @[Decode.scala 195:64]
  wire [3:0] imm_b_lo_hi_lo = io_inst[11:8]; // @[Decode.scala 195:78]
  wire [63:0] imm_b = {imm_b_hi_hi_hi,io_inst[31],imm_b_hi_lo,imm_b_lo_hi_hi,imm_b_lo_hi_lo,1'h0}; // @[Cat.scala 30:58]
  wire [31:0] imm_u_hi_hi = io_inst[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [19:0] imm_u_hi_lo = io_inst[31:12]; // @[Decode.scala 196:45]
  wire [63:0] imm_u = {imm_u_hi_hi,imm_u_hi_lo,12'h0}; // @[Cat.scala 30:58]
  wire [42:0] imm_j_hi_hi_hi = io_inst[31] ? 43'h7ffffffffff : 43'h0; // @[Bitwise.scala 72:12]
  wire [7:0] imm_j_hi_lo = io_inst[19:12]; // @[Decode.scala 197:55]
  wire  imm_j_lo_hi_hi = io_inst[20]; // @[Decode.scala 197:69]
  wire [9:0] imm_j_lo_hi_lo = io_inst[30:21]; // @[Decode.scala 197:79]
  wire [63:0] imm_j = {imm_j_hi_hi_hi,io_inst[31],imm_j_hi_lo,imm_j_lo_hi_hi,imm_j_lo_hi_lo,1'h0}; // @[Cat.scala 30:58]
  wire [63:0] _imm_T_3 = 6'h10 == inst_type ? imm_i : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _imm_T_5 = 6'h8 == inst_type ? imm_s : _imm_T_3; // @[Mux.scala 80:57]
  wire [63:0] _imm_T_7 = 6'h4 == inst_type ? imm_b : _imm_T_5; // @[Mux.scala 80:57]
  wire [63:0] _imm_T_9 = 6'h2 == inst_type ? imm_u : _imm_T_7; // @[Mux.scala 80:57]
  wire [63:0] imm = 6'h1 == inst_type ? imm_j : _imm_T_9; // @[Mux.scala 80:57]
  wire  _io_rs1_en_T = type_r | type_i; // @[Decode.scala 220:25]
  wire [63:0] _bu_jump_pc_T_2 = io_op1 + io_op2; // @[Decode.scala 232:59]
  wire [63:0] _bu_jump_pc_T_3 = _bu_jump_pc_T_2 & 64'hfffffffffffffffe; // @[Decode.scala 232:66]
  wire [63:0] _bu_jump_pc_T_5 = io_pc + imm; // @[Decode.scala 232:95]
  wire [63:0] bu_jump_pc = bu_code == 8'h80 ? _bu_jump_pc_T_3 : _bu_jump_pc_T_5; // @[Decode.scala 232:25]
  wire  _bu_jump_en_T = io_op1 == io_op2; // @[Decode.scala 234:31]
  wire  _bu_jump_en_T_1 = io_op1 != io_op2; // @[Decode.scala 235:31]
  wire  _bu_jump_en_T_4 = $signed(io_op1) < $signed(io_op2); // @[Decode.scala 236:41]
  wire  _bu_jump_en_T_7 = $signed(io_op1) >= $signed(io_op2); // @[Decode.scala 237:41]
  wire  _bu_jump_en_T_8 = io_op1 < io_op2; // @[Decode.scala 238:32]
  wire  _bu_jump_en_T_9 = io_op1 >= io_op2; // @[Decode.scala 239:32]
  wire  _bu_jump_en_T_13 = 8'h2 == bu_code ? _bu_jump_en_T_1 : 8'h1 == bu_code & _bu_jump_en_T; // @[Mux.scala 80:57]
  wire  _bu_jump_en_T_15 = 8'h4 == bu_code ? _bu_jump_en_T_4 : _bu_jump_en_T_13; // @[Mux.scala 80:57]
  wire  _bu_jump_en_T_17 = 8'h8 == bu_code ? _bu_jump_en_T_7 : _bu_jump_en_T_15; // @[Mux.scala 80:57]
  wire  _bu_jump_en_T_19 = 8'h10 == bu_code ? _bu_jump_en_T_8 : _bu_jump_en_T_17; // @[Mux.scala 80:57]
  wire  _bu_jump_en_T_21 = 8'h20 == bu_code ? _bu_jump_en_T_9 : _bu_jump_en_T_19; // @[Mux.scala 80:57]
  wire  bu_jump_en = 8'h80 == bu_code | (8'h40 == bu_code | _bu_jump_en_T_21); // @[Mux.scala 80:57]
  wire [63:0] _csru_jump_pc_T_1 = 7'h1 == csru_code ? io_mtvec : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] csru_jump_pc = 7'h2 == csru_code ? io_mepc : _csru_jump_pc_T_1; // @[Mux.scala 80:57]
  wire  csru_jump_en = 7'h2 == csru_code | 7'h1 == csru_code; // @[Mux.scala 80:57]
  assign io_rs1_en = type_r | type_i | type_s | type_b; // @[Decode.scala 220:45]
  assign io_rs2_en = type_r | type_s | type_b; // @[Decode.scala 221:35]
  assign io_rs1_addr = io_inst[19:15]; // @[Decode.scala 216:24]
  assign io_rs2_addr = io_inst[24:20]; // @[Decode.scala 217:24]
  assign io_rd_en = _io_rs1_en_T | type_u | jal; // @[Decode.scala 222:45]
  assign io_rd_addr = io_inst[11:7]; // @[Decode.scala 218:24]
  assign io_decode_info_fu_code = {fu_code_hi,fu_code_lo}; // @[Cat.scala 30:58]
  assign io_decode_info_alu_code = {alu_code_hi,alu_code_lo}; // @[Cat.scala 30:58]
  assign io_decode_info_bu_code = {bu_code_hi,bu_code_lo}; // @[Cat.scala 30:58]
  assign io_decode_info_lu_code = {lu_code_hi,lu_code_lo}; // @[Cat.scala 30:58]
  assign io_decode_info_su_code = {su_code_hi,su_code_lo}; // @[Cat.scala 30:58]
  assign io_decode_info_mdu_code = {mdu_code_hi,mdu_code_lo}; // @[Cat.scala 30:58]
  assign io_decode_info_csru_code = {csru_code_hi,csru_code_lo}; // @[Cat.scala 30:58]
  assign io_jump_en = bu_jump_en | csru_jump_en; // @[Decode.scala 253:30]
  assign io_jump_pc = bu_jump_en ? bu_jump_pc : csru_jump_pc; // @[Decode.scala 254:22]
  assign io_op1 = io_rs1_en ? io_rs1_data : 64'h0; // @[Decode.scala 224:18]
  assign io_op2 = io_rs2_en ? io_rs2_data : imm; // @[Decode.scala 225:18]
  assign io_imm = 6'h1 == inst_type ? imm_j : _imm_T_9; // @[Mux.scala 80:57]
  assign io_putch = io_inst == 32'h7b; // @[Decode.scala 124:24]
endmodule
module Execution(
  input  [15:0] io_decode_info_alu_code,
  input  [7:0]  io_decode_info_bu_code,
  input  [9:0]  io_decode_info_mdu_code,
  input  [6:0]  io_decode_info_csru_code,
  input  [63:0] io_op1,
  input  [63:0] io_op2,
  input  [63:0] io_pc,
  output [63:0] io_alu_out,
  output [63:0] io_bu_out,
  output [63:0] io_mdu_out,
  output [63:0] io_csru_out,
  input  [4:0]  io_rs1_addr,
  output [11:0] io_csr_raddr,
  input  [63:0] io_csr_rdata,
  output        io_csr_wen,
  output [11:0] io_csr_waddr,
  output [63:0] io_csr_wdata
);
  wire [63:0] _alu_out_T_1 = io_op1 + io_op2; // @[Execution.scala 51:39]
  wire [31:0] alu_out_hi = _alu_out_T_1[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] alu_out_lo = _alu_out_T_1[31:0]; // @[Execution.scala 41:41]
  wire [63:0] _alu_out_T_6 = {alu_out_hi,alu_out_lo}; // @[Cat.scala 30:58]
  wire [63:0] _alu_out_T_8 = io_op1 - io_op2; // @[Execution.scala 53:39]
  wire [31:0] alu_out_hi_1 = _alu_out_T_8[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] alu_out_lo_1 = _alu_out_T_8[31:0]; // @[Execution.scala 41:41]
  wire [63:0] _alu_out_T_13 = {alu_out_hi_1,alu_out_lo_1}; // @[Cat.scala 30:58]
  wire [63:0] _alu_out_T_15 = io_op2 + io_pc; // @[Execution.scala 55:39]
  wire [126:0] _GEN_0 = {{63'd0}, io_op1}; // @[Execution.scala 56:39]
  wire [126:0] _alu_out_T_17 = _GEN_0 << io_op2[5:0]; // @[Execution.scala 56:39]
  wire [63:0] _alu_out_T_20 = io_op1 >> io_op2[5:0]; // @[Execution.scala 57:39]
  wire [63:0] _alu_out_T_24 = $signed(io_op1) >>> io_op2[5:0]; // @[Execution.scala 58:68]
  wire [62:0] _GEN_1 = {{31'd0}, io_op1[31:0]}; // @[Execution.scala 59:51]
  wire [62:0] _alu_out_T_27 = _GEN_1 << io_op2[4:0]; // @[Execution.scala 59:51]
  wire [31:0] alu_out_hi_2 = _alu_out_T_27[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] alu_out_lo_2 = _alu_out_T_27[31:0]; // @[Execution.scala 41:41]
  wire [63:0] _alu_out_T_30 = {alu_out_hi_2,alu_out_lo_2}; // @[Cat.scala 30:58]
  wire [31:0] alu_out_lo_3 = io_op1[31:0] >> io_op2[4:0]; // @[Execution.scala 60:51]
  wire [31:0] alu_out_hi_3 = alu_out_lo_3[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _alu_out_T_36 = {alu_out_hi_3,alu_out_lo_3}; // @[Cat.scala 30:58]
  wire [31:0] _alu_out_T_38 = io_op1[31:0]; // @[Execution.scala 61:57]
  wire [31:0] alu_out_lo_4 = $signed(_alu_out_T_38) >>> io_op2[4:0]; // @[Execution.scala 61:80]
  wire [31:0] alu_out_hi_4 = alu_out_lo_4[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _alu_out_T_44 = {alu_out_hi_4,alu_out_lo_4}; // @[Cat.scala 30:58]
  wire [63:0] _alu_out_T_45 = io_op1 ^ io_op2; // @[Execution.scala 62:39]
  wire [63:0] _alu_out_T_46 = io_op1 | io_op2; // @[Execution.scala 63:39]
  wire [63:0] _alu_out_T_47 = io_op1 & io_op2; // @[Execution.scala 64:39]
  wire  _alu_out_T_50 = $signed(io_op1) < $signed(io_op2); // @[Execution.scala 65:48]
  wire  _alu_out_T_51 = io_op1 < io_op2; // @[Execution.scala 66:39]
  wire [63:0] _alu_out_T_53 = 16'h1 == io_decode_info_alu_code ? _alu_out_T_1 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _alu_out_T_55 = 16'h2 == io_decode_info_alu_code ? _alu_out_T_6 : _alu_out_T_53; // @[Mux.scala 80:57]
  wire [63:0] _alu_out_T_57 = 16'h4 == io_decode_info_alu_code ? _alu_out_T_8 : _alu_out_T_55; // @[Mux.scala 80:57]
  wire [63:0] _alu_out_T_59 = 16'h8 == io_decode_info_alu_code ? _alu_out_T_13 : _alu_out_T_57; // @[Mux.scala 80:57]
  wire [63:0] _alu_out_T_61 = 16'h10 == io_decode_info_alu_code ? _alu_out_T_15 : _alu_out_T_59; // @[Mux.scala 80:57]
  wire [63:0] _alu_out_T_63 = 16'h20 == io_decode_info_alu_code ? _alu_out_T_17[63:0] : _alu_out_T_61; // @[Mux.scala 80:57]
  wire [63:0] _alu_out_T_65 = 16'h40 == io_decode_info_alu_code ? _alu_out_T_20 : _alu_out_T_63; // @[Mux.scala 80:57]
  wire [63:0] _alu_out_T_67 = 16'h80 == io_decode_info_alu_code ? _alu_out_T_24 : _alu_out_T_65; // @[Mux.scala 80:57]
  wire [63:0] _alu_out_T_69 = 16'h100 == io_decode_info_alu_code ? _alu_out_T_30 : _alu_out_T_67; // @[Mux.scala 80:57]
  wire [63:0] _alu_out_T_71 = 16'h200 == io_decode_info_alu_code ? _alu_out_T_36 : _alu_out_T_69; // @[Mux.scala 80:57]
  wire [63:0] _alu_out_T_73 = 16'h400 == io_decode_info_alu_code ? _alu_out_T_44 : _alu_out_T_71; // @[Mux.scala 80:57]
  wire [63:0] _alu_out_T_75 = 16'h800 == io_decode_info_alu_code ? _alu_out_T_45 : _alu_out_T_73; // @[Mux.scala 80:57]
  wire [63:0] _alu_out_T_77 = 16'h1000 == io_decode_info_alu_code ? _alu_out_T_46 : _alu_out_T_75; // @[Mux.scala 80:57]
  wire [63:0] _alu_out_T_79 = 16'h2000 == io_decode_info_alu_code ? _alu_out_T_47 : _alu_out_T_77; // @[Mux.scala 80:57]
  wire [63:0] _alu_out_T_81 = 16'h4000 == io_decode_info_alu_code ? {{63'd0}, _alu_out_T_50} : _alu_out_T_79; // @[Mux.scala 80:57]
  wire [63:0] _bu_out_T_4 = io_pc + 64'h4; // @[Execution.scala 70:81]
  wire [127:0] _mdu_out_T = io_op1 * io_op2; // @[Execution.scala 74:33]
  wire [31:0] mdu_out_hi = _mdu_out_T[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] mdu_out_lo = _mdu_out_T[31:0]; // @[Execution.scala 41:41]
  wire [63:0] _mdu_out_T_4 = {mdu_out_hi,mdu_out_lo}; // @[Cat.scala 30:58]
  wire [64:0] _mdu_out_T_8 = $signed(io_op1) / $signed(io_op2); // @[Execution.scala 76:64]
  wire [31:0] _mdu_out_T_12 = io_op2[31:0]; // @[Execution.scala 77:68]
  wire [32:0] _mdu_out_T_14 = $signed(_alu_out_T_38) / $signed(_mdu_out_T_12); // @[Execution.scala 77:78]
  wire [63:0] _mdu_out_T_15 = io_op1 / io_op2; // @[Execution.scala 78:33]
  wire [31:0] _mdu_out_T_18 = io_op1[31:0] / io_op2[31:0]; // @[Execution.scala 79:40]
  wire [63:0] _mdu_out_T_22 = $signed(io_op1) % $signed(io_op2); // @[Execution.scala 80:64]
  wire [31:0] _mdu_out_T_28 = $signed(_alu_out_T_38) % $signed(_mdu_out_T_12); // @[Execution.scala 81:78]
  wire [63:0] _GEN_2 = io_op1 % io_op2; // @[Execution.scala 82:33]
  wire [63:0] _mdu_out_T_29 = _GEN_2[63:0]; // @[Execution.scala 82:33]
  wire [31:0] _GEN_3 = io_op1[31:0] % io_op2[31:0]; // @[Execution.scala 83:40]
  wire [31:0] _mdu_out_T_32 = _GEN_3[31:0]; // @[Execution.scala 83:40]
  wire [127:0] _mdu_out_T_34 = 10'h1 == io_decode_info_mdu_code ? _mdu_out_T : 128'h0; // @[Mux.scala 80:57]
  wire [127:0] _mdu_out_T_36 = 10'h2 == io_decode_info_mdu_code ? {{64'd0}, _mdu_out_T_4} : _mdu_out_T_34; // @[Mux.scala 80:57]
  wire [127:0] _mdu_out_T_38 = 10'h4 == io_decode_info_mdu_code ? {{63'd0}, _mdu_out_T_8} : _mdu_out_T_36; // @[Mux.scala 80:57]
  wire [127:0] _mdu_out_T_40 = 10'h8 == io_decode_info_mdu_code ? {{95'd0}, _mdu_out_T_14} : _mdu_out_T_38; // @[Mux.scala 80:57]
  wire [127:0] _mdu_out_T_42 = 10'h10 == io_decode_info_mdu_code ? {{64'd0}, _mdu_out_T_15} : _mdu_out_T_40; // @[Mux.scala 80:57]
  wire [127:0] _mdu_out_T_44 = 10'h20 == io_decode_info_mdu_code ? {{96'd0}, _mdu_out_T_18} : _mdu_out_T_42; // @[Mux.scala 80:57]
  wire [127:0] _mdu_out_T_46 = 10'h40 == io_decode_info_mdu_code ? {{64'd0}, _mdu_out_T_22} : _mdu_out_T_44; // @[Mux.scala 80:57]
  wire [127:0] _mdu_out_T_48 = 10'h80 == io_decode_info_mdu_code ? {{96'd0}, _mdu_out_T_28} : _mdu_out_T_46; // @[Mux.scala 80:57]
  wire [127:0] _mdu_out_T_50 = 10'h100 == io_decode_info_mdu_code ? {{64'd0}, _mdu_out_T_29} : _mdu_out_T_48; // @[Mux.scala 80:57]
  wire [127:0] mdu_out = 10'h200 == io_decode_info_mdu_code ? {{96'd0}, _mdu_out_T_32} : _mdu_out_T_50; // @[Mux.scala 80:57]
  wire [63:0] _csru_out_T_1 = 7'h4 == io_decode_info_csru_code ? io_csr_rdata : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _csru_out_T_3 = 7'h8 == io_decode_info_csru_code ? io_csr_rdata : _csru_out_T_1; // @[Mux.scala 80:57]
  wire [63:0] _csru_out_T_5 = 7'h10 == io_decode_info_csru_code ? io_csr_rdata : _csru_out_T_3; // @[Mux.scala 80:57]
  wire [63:0] _csru_out_T_7 = 7'h20 == io_decode_info_csru_code ? io_csr_rdata : _csru_out_T_5; // @[Mux.scala 80:57]
  wire [63:0] _csr_waddr_T_1 = 7'h4 == io_decode_info_csru_code ? io_op2 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _csr_waddr_T_3 = 7'h8 == io_decode_info_csru_code ? io_op2 : _csr_waddr_T_1; // @[Mux.scala 80:57]
  wire [63:0] _csr_waddr_T_5 = 7'h10 == io_decode_info_csru_code ? io_op2 : _csr_waddr_T_3; // @[Mux.scala 80:57]
  wire [63:0] _csr_waddr_T_7 = 7'h20 == io_decode_info_csru_code ? io_op2 : _csr_waddr_T_5; // @[Mux.scala 80:57]
  wire [63:0] csr_waddr = 7'h40 == io_decode_info_csru_code ? io_op2 : _csr_waddr_T_7; // @[Mux.scala 80:57]
  wire [63:0] _csr_wdata_T = io_csr_rdata | io_op1; // @[Execution.scala 110:39]
  wire [63:0] _csr_wdata_T_1 = ~io_op1; // @[Execution.scala 112:42]
  wire [63:0] _csr_wdata_T_2 = io_csr_rdata & _csr_wdata_T_1; // @[Execution.scala 112:39]
  wire [63:0] _csr_wdata_T_3 = {59'h0,io_rs1_addr}; // @[Cat.scala 30:58]
  wire [63:0] _csr_wdata_T_5 = ~_csr_wdata_T_3; // @[Execution.scala 114:42]
  wire [63:0] _csr_wdata_T_6 = io_csr_rdata & _csr_wdata_T_5; // @[Execution.scala 114:39]
  wire [63:0] _csr_wdata_T_8 = 7'h4 == io_decode_info_csru_code ? _csr_wdata_T : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _csr_wdata_T_10 = 7'h8 == io_decode_info_csru_code ? io_op1 : _csr_wdata_T_8; // @[Mux.scala 80:57]
  wire [63:0] _csr_wdata_T_12 = 7'h10 == io_decode_info_csru_code ? _csr_wdata_T_2 : _csr_wdata_T_10; // @[Mux.scala 80:57]
  wire [63:0] _csr_wdata_T_14 = 7'h20 == io_decode_info_csru_code ? _csr_wdata_T_3 : _csr_wdata_T_12; // @[Mux.scala 80:57]
  assign io_alu_out = 16'h8000 == io_decode_info_alu_code ? {{63'd0}, _alu_out_T_51} : _alu_out_T_81; // @[Mux.scala 80:57]
  assign io_bu_out = io_decode_info_bu_code == 8'h80 | io_decode_info_bu_code == 8'h40 ? _bu_out_T_4 : 64'h0; // @[Execution.scala 70:21]
  assign io_mdu_out = mdu_out[63:0]; // @[Execution.scala 120:17]
  assign io_csru_out = 7'h40 == io_decode_info_csru_code ? io_csr_rdata : _csru_out_T_7; // @[Mux.scala 80:57]
  assign io_csr_raddr = io_op2[11:0]; // @[Execution.scala 87:18]
  assign io_csr_wen = 7'h40 == io_decode_info_csru_code | (7'h20 == io_decode_info_csru_code | (7'h10 ==
    io_decode_info_csru_code | (7'h8 == io_decode_info_csru_code | 7'h4 == io_decode_info_csru_code))); // @[Mux.scala 80:57]
  assign io_csr_waddr = csr_waddr[11:0]; // @[Execution.scala 125:21]
  assign io_csr_wdata = 7'h40 == io_decode_info_csru_code ? _csr_wdata_T_6 : _csr_wdata_T_14; // @[Mux.scala 80:57]
endmodule
module RegFile(
  input         clock,
  input         reset,
  input  [4:0]  io_rs1_addr,
  input  [4:0]  io_rs2_addr,
  output [63:0] io_rs1_data,
  output [63:0] io_rs2_data,
  input  [4:0]  io_rd_addr,
  input  [63:0] io_rd_data,
  input         io_rd_en,
  output [63:0] rf_10
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  wire  dt_ar_clock; // @[RegFile.scala 25:21]
  wire [7:0] dt_ar_coreid; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_0; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_1; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_2; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_3; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_4; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_5; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_6; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_7; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_8; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_9; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_10; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_11; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_12; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_13; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_14; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_15; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_16; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_17; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_18; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_19; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_20; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_21; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_22; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_23; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_24; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_25; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_26; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_27; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_28; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_29; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_30; // @[RegFile.scala 25:21]
  wire [63:0] dt_ar_gpr_31; // @[RegFile.scala 25:21]
  reg [63:0] rf__0; // @[RegFile.scala 16:19]
  reg [63:0] rf__1; // @[RegFile.scala 16:19]
  reg [63:0] rf__2; // @[RegFile.scala 16:19]
  reg [63:0] rf__3; // @[RegFile.scala 16:19]
  reg [63:0] rf__4; // @[RegFile.scala 16:19]
  reg [63:0] rf__5; // @[RegFile.scala 16:19]
  reg [63:0] rf__6; // @[RegFile.scala 16:19]
  reg [63:0] rf__7; // @[RegFile.scala 16:19]
  reg [63:0] rf__8; // @[RegFile.scala 16:19]
  reg [63:0] rf__9; // @[RegFile.scala 16:19]
  reg [63:0] rf__10; // @[RegFile.scala 16:19]
  reg [63:0] rf__11; // @[RegFile.scala 16:19]
  reg [63:0] rf__12; // @[RegFile.scala 16:19]
  reg [63:0] rf__13; // @[RegFile.scala 16:19]
  reg [63:0] rf__14; // @[RegFile.scala 16:19]
  reg [63:0] rf__15; // @[RegFile.scala 16:19]
  reg [63:0] rf__16; // @[RegFile.scala 16:19]
  reg [63:0] rf__17; // @[RegFile.scala 16:19]
  reg [63:0] rf__18; // @[RegFile.scala 16:19]
  reg [63:0] rf__19; // @[RegFile.scala 16:19]
  reg [63:0] rf__20; // @[RegFile.scala 16:19]
  reg [63:0] rf__21; // @[RegFile.scala 16:19]
  reg [63:0] rf__22; // @[RegFile.scala 16:19]
  reg [63:0] rf__23; // @[RegFile.scala 16:19]
  reg [63:0] rf__24; // @[RegFile.scala 16:19]
  reg [63:0] rf__25; // @[RegFile.scala 16:19]
  reg [63:0] rf__26; // @[RegFile.scala 16:19]
  reg [63:0] rf__27; // @[RegFile.scala 16:19]
  reg [63:0] rf__28; // @[RegFile.scala 16:19]
  reg [63:0] rf__29; // @[RegFile.scala 16:19]
  reg [63:0] rf__30; // @[RegFile.scala 16:19]
  reg [63:0] rf__31; // @[RegFile.scala 16:19]
  wire [63:0] _GEN_65 = 5'h1 == io_rs1_addr ? rf__1 : rf__0; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_66 = 5'h2 == io_rs1_addr ? rf__2 : _GEN_65; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_67 = 5'h3 == io_rs1_addr ? rf__3 : _GEN_66; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_68 = 5'h4 == io_rs1_addr ? rf__4 : _GEN_67; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_69 = 5'h5 == io_rs1_addr ? rf__5 : _GEN_68; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_70 = 5'h6 == io_rs1_addr ? rf__6 : _GEN_69; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_71 = 5'h7 == io_rs1_addr ? rf__7 : _GEN_70; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_72 = 5'h8 == io_rs1_addr ? rf__8 : _GEN_71; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_73 = 5'h9 == io_rs1_addr ? rf__9 : _GEN_72; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_74 = 5'ha == io_rs1_addr ? rf__10 : _GEN_73; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_75 = 5'hb == io_rs1_addr ? rf__11 : _GEN_74; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_76 = 5'hc == io_rs1_addr ? rf__12 : _GEN_75; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_77 = 5'hd == io_rs1_addr ? rf__13 : _GEN_76; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_78 = 5'he == io_rs1_addr ? rf__14 : _GEN_77; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_79 = 5'hf == io_rs1_addr ? rf__15 : _GEN_78; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_80 = 5'h10 == io_rs1_addr ? rf__16 : _GEN_79; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_81 = 5'h11 == io_rs1_addr ? rf__17 : _GEN_80; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_82 = 5'h12 == io_rs1_addr ? rf__18 : _GEN_81; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_83 = 5'h13 == io_rs1_addr ? rf__19 : _GEN_82; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_84 = 5'h14 == io_rs1_addr ? rf__20 : _GEN_83; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_85 = 5'h15 == io_rs1_addr ? rf__21 : _GEN_84; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_86 = 5'h16 == io_rs1_addr ? rf__22 : _GEN_85; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_87 = 5'h17 == io_rs1_addr ? rf__23 : _GEN_86; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_88 = 5'h18 == io_rs1_addr ? rf__24 : _GEN_87; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_89 = 5'h19 == io_rs1_addr ? rf__25 : _GEN_88; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_90 = 5'h1a == io_rs1_addr ? rf__26 : _GEN_89; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_91 = 5'h1b == io_rs1_addr ? rf__27 : _GEN_90; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_92 = 5'h1c == io_rs1_addr ? rf__28 : _GEN_91; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_93 = 5'h1d == io_rs1_addr ? rf__29 : _GEN_92; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_94 = 5'h1e == io_rs1_addr ? rf__30 : _GEN_93; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_95 = 5'h1f == io_rs1_addr ? rf__31 : _GEN_94; // @[RegFile.scala 22:21 RegFile.scala 22:21]
  wire [63:0] _GEN_97 = 5'h1 == io_rs2_addr ? rf__1 : rf__0; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_98 = 5'h2 == io_rs2_addr ? rf__2 : _GEN_97; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_99 = 5'h3 == io_rs2_addr ? rf__3 : _GEN_98; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_100 = 5'h4 == io_rs2_addr ? rf__4 : _GEN_99; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_101 = 5'h5 == io_rs2_addr ? rf__5 : _GEN_100; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_102 = 5'h6 == io_rs2_addr ? rf__6 : _GEN_101; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_103 = 5'h7 == io_rs2_addr ? rf__7 : _GEN_102; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_104 = 5'h8 == io_rs2_addr ? rf__8 : _GEN_103; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_105 = 5'h9 == io_rs2_addr ? rf__9 : _GEN_104; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_106 = 5'ha == io_rs2_addr ? rf__10 : _GEN_105; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_107 = 5'hb == io_rs2_addr ? rf__11 : _GEN_106; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_108 = 5'hc == io_rs2_addr ? rf__12 : _GEN_107; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_109 = 5'hd == io_rs2_addr ? rf__13 : _GEN_108; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_110 = 5'he == io_rs2_addr ? rf__14 : _GEN_109; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_111 = 5'hf == io_rs2_addr ? rf__15 : _GEN_110; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_112 = 5'h10 == io_rs2_addr ? rf__16 : _GEN_111; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_113 = 5'h11 == io_rs2_addr ? rf__17 : _GEN_112; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_114 = 5'h12 == io_rs2_addr ? rf__18 : _GEN_113; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_115 = 5'h13 == io_rs2_addr ? rf__19 : _GEN_114; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_116 = 5'h14 == io_rs2_addr ? rf__20 : _GEN_115; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_117 = 5'h15 == io_rs2_addr ? rf__21 : _GEN_116; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_118 = 5'h16 == io_rs2_addr ? rf__22 : _GEN_117; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_119 = 5'h17 == io_rs2_addr ? rf__23 : _GEN_118; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_120 = 5'h18 == io_rs2_addr ? rf__24 : _GEN_119; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_121 = 5'h19 == io_rs2_addr ? rf__25 : _GEN_120; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_122 = 5'h1a == io_rs2_addr ? rf__26 : _GEN_121; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_123 = 5'h1b == io_rs2_addr ? rf__27 : _GEN_122; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_124 = 5'h1c == io_rs2_addr ? rf__28 : _GEN_123; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_125 = 5'h1d == io_rs2_addr ? rf__29 : _GEN_124; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_126 = 5'h1e == io_rs2_addr ? rf__30 : _GEN_125; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  wire [63:0] _GEN_127 = 5'h1f == io_rs2_addr ? rf__31 : _GEN_126; // @[RegFile.scala 23:21 RegFile.scala 23:21]
  DifftestArchIntRegState dt_ar ( // @[RegFile.scala 25:21]
    .clock(dt_ar_clock),
    .coreid(dt_ar_coreid),
    .gpr_0(dt_ar_gpr_0),
    .gpr_1(dt_ar_gpr_1),
    .gpr_2(dt_ar_gpr_2),
    .gpr_3(dt_ar_gpr_3),
    .gpr_4(dt_ar_gpr_4),
    .gpr_5(dt_ar_gpr_5),
    .gpr_6(dt_ar_gpr_6),
    .gpr_7(dt_ar_gpr_7),
    .gpr_8(dt_ar_gpr_8),
    .gpr_9(dt_ar_gpr_9),
    .gpr_10(dt_ar_gpr_10),
    .gpr_11(dt_ar_gpr_11),
    .gpr_12(dt_ar_gpr_12),
    .gpr_13(dt_ar_gpr_13),
    .gpr_14(dt_ar_gpr_14),
    .gpr_15(dt_ar_gpr_15),
    .gpr_16(dt_ar_gpr_16),
    .gpr_17(dt_ar_gpr_17),
    .gpr_18(dt_ar_gpr_18),
    .gpr_19(dt_ar_gpr_19),
    .gpr_20(dt_ar_gpr_20),
    .gpr_21(dt_ar_gpr_21),
    .gpr_22(dt_ar_gpr_22),
    .gpr_23(dt_ar_gpr_23),
    .gpr_24(dt_ar_gpr_24),
    .gpr_25(dt_ar_gpr_25),
    .gpr_26(dt_ar_gpr_26),
    .gpr_27(dt_ar_gpr_27),
    .gpr_28(dt_ar_gpr_28),
    .gpr_29(dt_ar_gpr_29),
    .gpr_30(dt_ar_gpr_30),
    .gpr_31(dt_ar_gpr_31)
  );
  assign io_rs1_data = io_rs1_addr != 5'h0 ? _GEN_95 : 64'h0; // @[RegFile.scala 22:21]
  assign io_rs2_data = io_rs2_addr != 5'h0 ? _GEN_127 : 64'h0; // @[RegFile.scala 23:21]
  assign rf_10 = rf__10;
  assign dt_ar_clock = clock; // @[RegFile.scala 26:19]
  assign dt_ar_coreid = 8'h0; // @[RegFile.scala 27:19]
  assign dt_ar_gpr_0 = rf__0; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_1 = rf__1; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_2 = rf__2; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_3 = rf__3; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_4 = rf__4; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_5 = rf__5; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_6 = rf__6; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_7 = rf__7; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_8 = rf__8; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_9 = rf__9; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_10 = rf__10; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_11 = rf__11; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_12 = rf__12; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_13 = rf__13; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_14 = rf__14; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_15 = rf__15; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_16 = rf__16; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_17 = rf__17; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_18 = rf__18; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_19 = rf__19; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_20 = rf__20; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_21 = rf__21; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_22 = rf__22; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_23 = rf__23; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_24 = rf__24; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_25 = rf__25; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_26 = rf__26; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_27 = rf__27; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_28 = rf__28; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_29 = rf__29; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_30 = rf__30; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_31 = rf__31; // @[RegFile.scala 28:19]
  always @(posedge clock) begin
    if (reset) begin // @[RegFile.scala 16:19]
      rf__0 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h0 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__0 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__1 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h1 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__1 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__2 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h2 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__2 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__3 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h3 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__3 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__4 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h4 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__4 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__5 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h5 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__5 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__6 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h6 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__6 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__7 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h7 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__7 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__8 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h8 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__8 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__9 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h9 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__9 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__10 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'ha == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__10 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__11 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'hb == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__11 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__12 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'hc == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__12 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__13 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'hd == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__13 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__14 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'he == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__14 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__15 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'hf == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__15 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__16 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h10 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__16 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__17 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h11 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__17 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__18 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h12 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__18 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__19 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h13 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__19 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__20 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h14 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__20 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__21 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h15 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__21 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__22 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h16 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__22 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__23 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h17 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__23 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__24 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h18 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__24 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__25 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h19 == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__25 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__26 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h1a == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__26 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__27 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h1b == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__27 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__28 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h1c == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__28 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__29 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h1d == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__29 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__30 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h1e == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__30 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
    if (reset) begin // @[RegFile.scala 16:19]
      rf__31 <= 64'h0; // @[RegFile.scala 16:19]
    end else if (io_rd_en & io_rd_addr != 5'h0) begin // @[RegFile.scala 18:43]
      if (5'h1f == io_rd_addr) begin // @[RegFile.scala 19:20]
        rf__31 <= io_rd_data; // @[RegFile.scala 19:20]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  rf__0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  rf__1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  rf__2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  rf__3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  rf__4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  rf__5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  rf__6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  rf__7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  rf__8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  rf__9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  rf__10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  rf__11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  rf__12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  rf__13 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  rf__14 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  rf__15 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  rf__16 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  rf__17 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  rf__18 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  rf__19 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  rf__20 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  rf__21 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  rf__22 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  rf__23 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  rf__24 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  rf__25 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  rf__26 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  rf__27 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  rf__28 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  rf__29 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  rf__30 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  rf__31 = _RAND_31[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Csr(
  input         clock,
  input         reset,
  input  [11:0] io_raddr,
  output [63:0] io_rdata,
  input         io_wen,
  input  [11:0] io_waddr,
  input  [63:0] io_wdata,
  input         io_csru_code_valid,
  input  [6:0]  io_csru_code,
  input  [63:0] io_pc,
  output [63:0] io_mtvec,
  output [63:0] io_mepc
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire  dt_cs_clock; // @[Csr.scala 100:23]
  wire [7:0] dt_cs_coreid; // @[Csr.scala 100:23]
  wire [1:0] dt_cs_priviledgeMode; // @[Csr.scala 100:23]
  wire [63:0] dt_cs_mstatus; // @[Csr.scala 100:23]
  wire [63:0] dt_cs_sstatus; // @[Csr.scala 100:23]
  wire [63:0] dt_cs_mepc; // @[Csr.scala 100:23]
  wire [63:0] dt_cs_sepc; // @[Csr.scala 100:23]
  wire [63:0] dt_cs_mtval; // @[Csr.scala 100:23]
  wire [63:0] dt_cs_stval; // @[Csr.scala 100:23]
  wire [63:0] dt_cs_mtvec; // @[Csr.scala 100:23]
  wire [63:0] dt_cs_stvec; // @[Csr.scala 100:23]
  wire [63:0] dt_cs_mcause; // @[Csr.scala 100:23]
  wire [63:0] dt_cs_scause; // @[Csr.scala 100:23]
  wire [63:0] dt_cs_satp; // @[Csr.scala 100:23]
  wire [63:0] dt_cs_mip; // @[Csr.scala 100:23]
  wire [63:0] dt_cs_mie; // @[Csr.scala 100:23]
  wire [63:0] dt_cs_mscratch; // @[Csr.scala 100:23]
  wire [63:0] dt_cs_sscratch; // @[Csr.scala 100:23]
  wire [63:0] dt_cs_mideleg; // @[Csr.scala 100:23]
  wire [63:0] dt_cs_medeleg; // @[Csr.scala 100:23]
  reg [63:0] mstatus; // @[Csr.scala 40:30]
  reg [63:0] mtvec; // @[Csr.scala 41:30]
  reg [63:0] mepc; // @[Csr.scala 42:30]
  reg [63:0] mcause; // @[Csr.scala 43:30]
  reg [63:0] mcycle; // @[Csr.scala 44:30]
  reg [63:0] mie; // @[Csr.scala 47:30]
  reg [63:0] mip; // @[Csr.scala 48:30]
  reg [63:0] mscratch; // @[Csr.scala 49:30]
  reg [63:0] satp; // @[Csr.scala 50:30]
  wire [63:0] _io_rdata_T_1 = 12'h300 == io_raddr ? mstatus : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _io_rdata_T_3 = 12'h305 == io_raddr ? mtvec : _io_rdata_T_1; // @[Mux.scala 80:57]
  wire [63:0] _io_rdata_T_5 = 12'h341 == io_raddr ? mepc : _io_rdata_T_3; // @[Mux.scala 80:57]
  wire [63:0] _io_rdata_T_7 = 12'h342 == io_raddr ? mcause : _io_rdata_T_5; // @[Mux.scala 80:57]
  wire [63:0] _mcycle_T_3 = mcycle + 64'h1; // @[Csr.scala 60:68]
  wire  mstatus_SD = io_wdata[14:13] == 2'h3 | io_wdata[16:15] == 2'h3; // @[Csr.scala 62:60]
  wire [62:0] mstatus_lo = io_wdata[62:0]; // @[Csr.scala 64:44]
  wire [63:0] _mstatus_T = {mstatus_SD,mstatus_lo}; // @[Cat.scala 30:58]
  wire  _T_3 = io_csru_code_valid & io_csru_code == 7'h1; // @[Csr.scala 66:34]
  wire [50:0] mstatus_hi_hi_hi = mstatus[63:13]; // @[Csr.scala 67:31]
  wire [2:0] mstatus_hi_lo_hi = mstatus[10:8]; // @[Csr.scala 67:61]
  wire  mstatus_hi_lo_lo = mstatus[3]; // @[Csr.scala 67:76]
  wire [2:0] mstatus_lo_hi_hi = mstatus[6:4]; // @[Csr.scala 67:88]
  wire [2:0] mstatus_lo_lo = mstatus[2:0]; // @[Csr.scala 67:108]
  wire [63:0] _mstatus_T_1 = {mstatus_hi_hi_hi,2'h3,mstatus_hi_lo_hi,mstatus_hi_lo_lo,mstatus_lo_hi_hi,1'h0,
    mstatus_lo_lo}; // @[Cat.scala 30:58]
  wire  mstatus_lo_hi_lo = mstatus[7]; // @[Csr.scala 70:96]
  wire [63:0] _mstatus_T_2 = {mstatus_hi_hi_hi,2'h0,mstatus_hi_lo_hi,1'h1,mstatus_lo_hi_hi,mstatus_lo_hi_lo,
    mstatus_lo_lo}; // @[Cat.scala 30:58]
  wire  _mcause_T_1 = io_wen & io_waddr == 12'h342; // @[Csr.scala 82:27]
  DifftestCSRState dt_cs ( // @[Csr.scala 100:23]
    .clock(dt_cs_clock),
    .coreid(dt_cs_coreid),
    .priviledgeMode(dt_cs_priviledgeMode),
    .mstatus(dt_cs_mstatus),
    .sstatus(dt_cs_sstatus),
    .mepc(dt_cs_mepc),
    .sepc(dt_cs_sepc),
    .mtval(dt_cs_mtval),
    .stval(dt_cs_stval),
    .mtvec(dt_cs_mtvec),
    .stvec(dt_cs_stvec),
    .mcause(dt_cs_mcause),
    .scause(dt_cs_scause),
    .satp(dt_cs_satp),
    .mip(dt_cs_mip),
    .mie(dt_cs_mie),
    .mscratch(dt_cs_mscratch),
    .sscratch(dt_cs_sscratch),
    .mideleg(dt_cs_mideleg),
    .medeleg(dt_cs_medeleg)
  );
  assign io_rdata = 12'hb00 == io_raddr ? mcycle : _io_rdata_T_7; // @[Mux.scala 80:57]
  assign io_mtvec = mtvec; // @[Csr.scala 94:14]
  assign io_mepc = mepc; // @[Csr.scala 95:14]
  assign dt_cs_clock = clock; // @[Csr.scala 101:29]
  assign dt_cs_coreid = 8'h0; // @[Csr.scala 102:29]
  assign dt_cs_priviledgeMode = 2'h3; // @[Csr.scala 103:29]
  assign dt_cs_mstatus = mstatus; // @[Csr.scala 104:29]
  assign dt_cs_sstatus = mstatus & 64'h80000003000de122; // @[Csr.scala 105:40]
  assign dt_cs_mepc = mepc; // @[Csr.scala 106:29]
  assign dt_cs_sepc = 64'h0; // @[Csr.scala 107:29]
  assign dt_cs_mtval = 64'h0; // @[Csr.scala 108:29]
  assign dt_cs_stval = 64'h0; // @[Csr.scala 109:29]
  assign dt_cs_mtvec = mtvec; // @[Csr.scala 110:29]
  assign dt_cs_stvec = 64'h0; // @[Csr.scala 111:29]
  assign dt_cs_mcause = mcause; // @[Csr.scala 112:29]
  assign dt_cs_scause = 64'h0; // @[Csr.scala 113:29]
  assign dt_cs_satp = satp; // @[Csr.scala 114:29]
  assign dt_cs_mip = mip; // @[Csr.scala 115:29]
  assign dt_cs_mie = mie; // @[Csr.scala 116:29]
  assign dt_cs_mscratch = mscratch; // @[Csr.scala 117:29]
  assign dt_cs_sscratch = 64'h0; // @[Csr.scala 118:29]
  assign dt_cs_mideleg = 64'h0; // @[Csr.scala 119:29]
  assign dt_cs_medeleg = 64'h0; // @[Csr.scala 120:29]
  always @(posedge clock) begin
    if (reset) begin // @[Csr.scala 40:30]
      mstatus <= 64'h1800; // @[Csr.scala 40:30]
    end else if (io_wen & io_waddr == 12'h300) begin // @[Csr.scala 63:41]
      mstatus <= _mstatus_T; // @[Csr.scala 64:17]
    end else if (io_csru_code_valid & io_csru_code == 7'h1) begin // @[Csr.scala 66:64]
      mstatus <= _mstatus_T_1; // @[Csr.scala 67:17]
    end else if (io_csru_code_valid & io_csru_code == 7'h2) begin // @[Csr.scala 69:64]
      mstatus <= _mstatus_T_2; // @[Csr.scala 70:17]
    end
    if (reset) begin // @[Csr.scala 41:30]
      mtvec <= 64'h0; // @[Csr.scala 41:30]
    end else if (io_wen & io_waddr == 12'h305) begin // @[Csr.scala 76:19]
      mtvec <= io_wdata;
    end
    if (reset) begin // @[Csr.scala 42:30]
      mepc <= 64'h0; // @[Csr.scala 42:30]
    end else if (io_wen & io_waddr == 12'h341) begin // @[Csr.scala 78:39]
      mepc <= io_wdata; // @[Csr.scala 78:45]
    end else if (_T_3) begin // @[Csr.scala 79:65]
      mepc <= io_pc; // @[Csr.scala 79:71]
    end
    if (reset) begin // @[Csr.scala 43:30]
      mcause <= 64'h0; // @[Csr.scala 43:30]
    end else if (_mcause_T_1) begin // @[Csr.scala 83:41]
      mcause <= io_wdata; // @[Csr.scala 83:49]
    end else if (_T_3) begin // @[Csr.scala 84:65]
      mcause <= 64'hb; // @[Csr.scala 84:73]
    end
    if (reset) begin // @[Csr.scala 44:30]
      mcycle <= 64'h0; // @[Csr.scala 44:30]
    end else if (io_wen & io_waddr == 12'hb00) begin // @[Csr.scala 60:19]
      mcycle <= io_wdata;
    end else begin
      mcycle <= _mcycle_T_3;
    end
    if (reset) begin // @[Csr.scala 47:30]
      mie <= 64'h0; // @[Csr.scala 47:30]
    end else if (io_wen & io_waddr == 12'h304) begin // @[Csr.scala 88:23]
      mie <= io_wdata;
    end
    if (reset) begin // @[Csr.scala 48:30]
      mip <= 64'h0; // @[Csr.scala 48:30]
    end else if (io_wen & io_waddr == 12'h344) begin // @[Csr.scala 89:23]
      mip <= io_wdata;
    end
    if (reset) begin // @[Csr.scala 49:30]
      mscratch <= 64'h0; // @[Csr.scala 49:30]
    end else if (io_wen & io_waddr == 12'h340) begin // @[Csr.scala 90:23]
      mscratch <= io_wdata;
    end
    if (reset) begin // @[Csr.scala 50:30]
      satp <= 64'h0; // @[Csr.scala 50:30]
    end else if (io_wen & io_waddr == 12'h180) begin // @[Csr.scala 91:23]
      satp <= io_wdata;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mstatus = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  mtvec = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  mepc = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  mcause = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  mcycle = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  mie = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  mip = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  mscratch = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  satp = _RAND_8[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PreAccessMemory(
  input  [6:0]  io_lu_code,
  input  [3:0]  io_su_code,
  input  [63:0] io_op1,
  input  [63:0] io_op2,
  input  [63:0] io_imm,
  output [5:0]  io_lu_shift,
  output        io_ren,
  output [63:0] io_raddr,
  output        io_wen,
  output [63:0] io_waddr,
  output [63:0] io_wdata,
  output [7:0]  io_wmask
);
  wire [63:0] lu_offset = io_op1 + io_op2; // @[PreAccessMemory.scala 23:28]
  wire [63:0] su_offset = io_op1 + io_imm; // @[PreAccessMemory.scala 29:28]
  wire [5:0] su_shift = {su_offset[2:0], 3'h0}; // @[PreAccessMemory.scala 30:37]
  wire [126:0] _GEN_0 = {{63'd0}, io_op2}; // @[PreAccessMemory.scala 33:28]
  wire [126:0] su_wdata = _GEN_0 << su_shift; // @[PreAccessMemory.scala 33:28]
  wire [7:0] _su_wmask_T_1 = 8'h1 << su_offset[2:0]; // @[PreAccessMemory.scala 35:37]
  wire [8:0] _su_wmask_T_3 = 9'h3 << su_offset[2:0]; // @[PreAccessMemory.scala 36:37]
  wire [10:0] _su_wmask_T_5 = 11'hf << su_offset[2:0]; // @[PreAccessMemory.scala 37:37]
  wire [7:0] _su_wmask_T_7 = 4'h1 == io_su_code ? _su_wmask_T_1 : 8'h0; // @[Mux.scala 80:57]
  wire [8:0] _su_wmask_T_9 = 4'h2 == io_su_code ? _su_wmask_T_3 : {{1'd0}, _su_wmask_T_7}; // @[Mux.scala 80:57]
  wire [10:0] _su_wmask_T_11 = 4'h4 == io_su_code ? _su_wmask_T_5 : {{2'd0}, _su_wmask_T_9}; // @[Mux.scala 80:57]
  wire [10:0] su_wmask = 4'h8 == io_su_code ? 11'hff : _su_wmask_T_11; // @[Mux.scala 80:57]
  assign io_lu_shift = {lu_offset[2:0], 3'h0}; // @[PreAccessMemory.scala 24:36]
  assign io_ren = io_lu_code != 7'h0; // @[PreAccessMemory.scala 25:29]
  assign io_raddr = lu_offset & 64'hfffffffffffffff8; // @[PreAccessMemory.scala 26:30]
  assign io_wen = io_su_code != 4'h0; // @[PreAccessMemory.scala 31:32]
  assign io_waddr = su_offset & 64'hfffffffffffffff8; // @[PreAccessMemory.scala 32:31]
  assign io_wdata = su_wdata[63:0]; // @[PreAccessMemory.scala 46:17]
  assign io_wmask = su_wmask[7:0]; // @[PreAccessMemory.scala 47:17]
endmodule
module AccessMemory(
  input  [6:0]  io_lu_code,
  input  [5:0]  io_lu_shift,
  input  [63:0] io_rdata,
  output [63:0] io_lu_out
);
  wire [63:0] _io_lu_out_T = io_rdata >> io_lu_shift; // @[AccessMemory.scala 23:41]
  wire [55:0] io_lu_out_hi = _io_lu_out_T[7] ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 72:12]
  wire [7:0] io_lu_out_lo = _io_lu_out_T[7:0]; // @[AccessMemory.scala 13:40]
  wire [63:0] _io_lu_out_T_3 = {io_lu_out_hi,io_lu_out_lo}; // @[Cat.scala 30:58]
  wire [47:0] io_lu_out_hi_1 = _io_lu_out_T[15] ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 72:12]
  wire [15:0] io_lu_out_lo_1 = _io_lu_out_T[15:0]; // @[AccessMemory.scala 14:41]
  wire [63:0] _io_lu_out_T_7 = {io_lu_out_hi_1,io_lu_out_lo_1}; // @[Cat.scala 30:58]
  wire [31:0] io_lu_out_hi_2 = _io_lu_out_T[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] io_lu_out_lo_2 = _io_lu_out_T[31:0]; // @[AccessMemory.scala 15:41]
  wire [63:0] _io_lu_out_T_11 = {io_lu_out_hi_2,io_lu_out_lo_2}; // @[Cat.scala 30:58]
  wire [63:0] _io_lu_out_T_14 = {56'h0,io_lu_out_lo}; // @[Cat.scala 30:58]
  wire [63:0] _io_lu_out_T_16 = {48'h0,io_lu_out_lo_1}; // @[Cat.scala 30:58]
  wire [63:0] _io_lu_out_T_18 = {32'h0,io_lu_out_lo_2}; // @[Cat.scala 30:58]
  wire [63:0] _io_lu_out_T_20 = 7'h1 == io_lu_code ? _io_lu_out_T_3 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _io_lu_out_T_22 = 7'h2 == io_lu_code ? _io_lu_out_T_7 : _io_lu_out_T_20; // @[Mux.scala 80:57]
  wire [63:0] _io_lu_out_T_24 = 7'h4 == io_lu_code ? _io_lu_out_T_11 : _io_lu_out_T_22; // @[Mux.scala 80:57]
  wire [63:0] _io_lu_out_T_26 = 7'h8 == io_lu_code ? _io_lu_out_T : _io_lu_out_T_24; // @[Mux.scala 80:57]
  wire [63:0] _io_lu_out_T_28 = 7'h10 == io_lu_code ? _io_lu_out_T_14 : _io_lu_out_T_26; // @[Mux.scala 80:57]
  wire [63:0] _io_lu_out_T_30 = 7'h20 == io_lu_code ? _io_lu_out_T_16 : _io_lu_out_T_28; // @[Mux.scala 80:57]
  assign io_lu_out = 7'h40 == io_lu_code ? _io_lu_out_T_18 : _io_lu_out_T_30; // @[Mux.scala 80:57]
endmodule
module WriteBack(
  input  [5:0]  io_fu_code,
  input  [63:0] io_alu_out,
  input  [63:0] io_bu_out,
  input  [63:0] io_mdu_out,
  input  [63:0] io_lu_out,
  input  [63:0] io_csru_out,
  output [63:0] io_out
);
  wire [63:0] _io_out_T_1 = 6'h1 == io_fu_code ? io_alu_out : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _io_out_T_3 = 6'h2 == io_fu_code ? io_bu_out : _io_out_T_1; // @[Mux.scala 80:57]
  wire [63:0] _io_out_T_5 = 6'h4 == io_fu_code ? io_lu_out : _io_out_T_3; // @[Mux.scala 80:57]
  wire [63:0] _io_out_T_7 = 6'h8 == io_fu_code ? 64'h0 : _io_out_T_5; // @[Mux.scala 80:57]
  wire [63:0] _io_out_T_9 = 6'h10 == io_fu_code ? io_mdu_out : _io_out_T_7; // @[Mux.scala 80:57]
  assign io_out = 6'h20 == io_fu_code ? io_csru_out : _io_out_T_9; // @[Mux.scala 80:57]
endmodule
module CorrelationConflict(
  input        io_rs_valid,
  input        io_rd_valid,
  input        io_rs1_en,
  input        io_rs2_en,
  input  [4:0] io_rs1_addr,
  input  [4:0] io_rs2_addr,
  input        io_rd_en,
  input  [4:0] io_rd_addr,
  output       io_conflict
);
  wire  inst_valid = io_rs_valid & io_rd_valid; // @[PipelineReg.scala 294:39]
  wire  rs1_conflict = io_rs1_en & io_rs1_addr == io_rd_addr; // @[PipelineReg.scala 295:37]
  wire  rs2_conflict = io_rs2_en & io_rs2_addr == io_rd_addr; // @[PipelineReg.scala 296:37]
  wire  rd_valid = io_rd_addr != 5'h0 & io_rd_en; // @[PipelineReg.scala 297:48]
  assign io_conflict = inst_valid & rd_valid & (rs1_conflict | rs2_conflict); // @[PipelineReg.scala 299:43]
endmodule
module RegfileConflict(
  input        io_rs_valid,
  input        io_rs1_en,
  input        io_rs2_en,
  input  [4:0] io_rs1_addr,
  input  [4:0] io_rs2_addr,
  input        io_rd1_valid,
  input        io_rd1_en,
  input  [4:0] io_rd1_addr,
  input        io_rd2_valid,
  input        io_rd2_en,
  input  [4:0] io_rd2_addr,
  input        io_rd3_valid,
  input        io_rd3_en,
  input  [4:0] io_rd3_addr,
  output       io_conflict
);
  wire  cconflict1_io_rs_valid; // @[PipelineReg.scala 322:28]
  wire  cconflict1_io_rd_valid; // @[PipelineReg.scala 322:28]
  wire  cconflict1_io_rs1_en; // @[PipelineReg.scala 322:28]
  wire  cconflict1_io_rs2_en; // @[PipelineReg.scala 322:28]
  wire [4:0] cconflict1_io_rs1_addr; // @[PipelineReg.scala 322:28]
  wire [4:0] cconflict1_io_rs2_addr; // @[PipelineReg.scala 322:28]
  wire  cconflict1_io_rd_en; // @[PipelineReg.scala 322:28]
  wire [4:0] cconflict1_io_rd_addr; // @[PipelineReg.scala 322:28]
  wire  cconflict1_io_conflict; // @[PipelineReg.scala 322:28]
  wire  cconflict2_io_rs_valid; // @[PipelineReg.scala 323:28]
  wire  cconflict2_io_rd_valid; // @[PipelineReg.scala 323:28]
  wire  cconflict2_io_rs1_en; // @[PipelineReg.scala 323:28]
  wire  cconflict2_io_rs2_en; // @[PipelineReg.scala 323:28]
  wire [4:0] cconflict2_io_rs1_addr; // @[PipelineReg.scala 323:28]
  wire [4:0] cconflict2_io_rs2_addr; // @[PipelineReg.scala 323:28]
  wire  cconflict2_io_rd_en; // @[PipelineReg.scala 323:28]
  wire [4:0] cconflict2_io_rd_addr; // @[PipelineReg.scala 323:28]
  wire  cconflict2_io_conflict; // @[PipelineReg.scala 323:28]
  wire  cconflict3_io_rs_valid; // @[PipelineReg.scala 324:28]
  wire  cconflict3_io_rd_valid; // @[PipelineReg.scala 324:28]
  wire  cconflict3_io_rs1_en; // @[PipelineReg.scala 324:28]
  wire  cconflict3_io_rs2_en; // @[PipelineReg.scala 324:28]
  wire [4:0] cconflict3_io_rs1_addr; // @[PipelineReg.scala 324:28]
  wire [4:0] cconflict3_io_rs2_addr; // @[PipelineReg.scala 324:28]
  wire  cconflict3_io_rd_en; // @[PipelineReg.scala 324:28]
  wire [4:0] cconflict3_io_rd_addr; // @[PipelineReg.scala 324:28]
  wire  cconflict3_io_conflict; // @[PipelineReg.scala 324:28]
  CorrelationConflict cconflict1 ( // @[PipelineReg.scala 322:28]
    .io_rs_valid(cconflict1_io_rs_valid),
    .io_rd_valid(cconflict1_io_rd_valid),
    .io_rs1_en(cconflict1_io_rs1_en),
    .io_rs2_en(cconflict1_io_rs2_en),
    .io_rs1_addr(cconflict1_io_rs1_addr),
    .io_rs2_addr(cconflict1_io_rs2_addr),
    .io_rd_en(cconflict1_io_rd_en),
    .io_rd_addr(cconflict1_io_rd_addr),
    .io_conflict(cconflict1_io_conflict)
  );
  CorrelationConflict cconflict2 ( // @[PipelineReg.scala 323:28]
    .io_rs_valid(cconflict2_io_rs_valid),
    .io_rd_valid(cconflict2_io_rd_valid),
    .io_rs1_en(cconflict2_io_rs1_en),
    .io_rs2_en(cconflict2_io_rs2_en),
    .io_rs1_addr(cconflict2_io_rs1_addr),
    .io_rs2_addr(cconflict2_io_rs2_addr),
    .io_rd_en(cconflict2_io_rd_en),
    .io_rd_addr(cconflict2_io_rd_addr),
    .io_conflict(cconflict2_io_conflict)
  );
  CorrelationConflict cconflict3 ( // @[PipelineReg.scala 324:28]
    .io_rs_valid(cconflict3_io_rs_valid),
    .io_rd_valid(cconflict3_io_rd_valid),
    .io_rs1_en(cconflict3_io_rs1_en),
    .io_rs2_en(cconflict3_io_rs2_en),
    .io_rs1_addr(cconflict3_io_rs1_addr),
    .io_rs2_addr(cconflict3_io_rs2_addr),
    .io_rd_en(cconflict3_io_rd_en),
    .io_rd_addr(cconflict3_io_rd_addr),
    .io_conflict(cconflict3_io_conflict)
  );
  assign io_conflict = cconflict1_io_conflict | cconflict2_io_conflict | cconflict3_io_conflict; // @[PipelineReg.scala 353:69]
  assign cconflict1_io_rs_valid = io_rs_valid; // @[PipelineReg.scala 326:29]
  assign cconflict1_io_rd_valid = io_rd1_valid; // @[PipelineReg.scala 327:29]
  assign cconflict1_io_rs1_en = io_rs1_en; // @[PipelineReg.scala 328:29]
  assign cconflict1_io_rs2_en = io_rs2_en; // @[PipelineReg.scala 329:29]
  assign cconflict1_io_rs1_addr = io_rs1_addr; // @[PipelineReg.scala 330:29]
  assign cconflict1_io_rs2_addr = io_rs2_addr; // @[PipelineReg.scala 331:29]
  assign cconflict1_io_rd_en = io_rd1_en; // @[PipelineReg.scala 332:29]
  assign cconflict1_io_rd_addr = io_rd1_addr; // @[PipelineReg.scala 333:29]
  assign cconflict2_io_rs_valid = io_rs_valid; // @[PipelineReg.scala 335:29]
  assign cconflict2_io_rd_valid = io_rd2_valid; // @[PipelineReg.scala 336:29]
  assign cconflict2_io_rs1_en = io_rs1_en; // @[PipelineReg.scala 337:29]
  assign cconflict2_io_rs2_en = io_rs2_en; // @[PipelineReg.scala 338:29]
  assign cconflict2_io_rs1_addr = io_rs1_addr; // @[PipelineReg.scala 339:29]
  assign cconflict2_io_rs2_addr = io_rs2_addr; // @[PipelineReg.scala 340:29]
  assign cconflict2_io_rd_en = io_rd2_en; // @[PipelineReg.scala 341:29]
  assign cconflict2_io_rd_addr = io_rd2_addr; // @[PipelineReg.scala 342:29]
  assign cconflict3_io_rs_valid = io_rs_valid; // @[PipelineReg.scala 344:29]
  assign cconflict3_io_rd_valid = io_rd3_valid; // @[PipelineReg.scala 345:29]
  assign cconflict3_io_rs1_en = io_rs1_en; // @[PipelineReg.scala 346:29]
  assign cconflict3_io_rs2_en = io_rs2_en; // @[PipelineReg.scala 347:29]
  assign cconflict3_io_rs1_addr = io_rs1_addr; // @[PipelineReg.scala 348:29]
  assign cconflict3_io_rs2_addr = io_rs2_addr; // @[PipelineReg.scala 349:29]
  assign cconflict3_io_rd_en = io_rd3_en; // @[PipelineReg.scala 350:29]
  assign cconflict3_io_rd_addr = io_rd3_addr; // @[PipelineReg.scala 351:29]
endmodule
module ImemoryReadHold(
  input         clock,
  input         reset,
  input         io_ren,
  input  [63:0] io_raddr,
  output [63:0] io_imem_raddr
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] raddr; // @[Reg.scala 27:20]
  assign io_imem_raddr = io_ren ? io_raddr : raddr; // @[PipelineReg.scala 276:23]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 27:20]
      raddr <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_ren) begin // @[Reg.scala 28:19]
      raddr <= io_raddr; // @[Reg.scala 28:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  raddr = _RAND_0[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IDReg(
  input         clock,
  input         reset,
  output [63:0] io_imem_addr,
  input  [31:0] io_imem_data,
  input         io_pr_valid_in,
  output        io_pr_valid_out,
  input         io_pr_en,
  input  [63:0] io_pc_in,
  output [63:0] io_pc_out,
  output [31:0] io_inst_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  imemrh_clock; // @[PipelineReg.scala 23:25]
  wire  imemrh_reset; // @[PipelineReg.scala 23:25]
  wire  imemrh_io_ren; // @[PipelineReg.scala 23:25]
  wire [63:0] imemrh_io_raddr; // @[PipelineReg.scala 23:25]
  wire [63:0] imemrh_io_imem_raddr; // @[PipelineReg.scala 23:25]
  reg  valid; // @[Reg.scala 27:20]
  reg [63:0] pc; // @[Reg.scala 27:20]
  ImemoryReadHold imemrh ( // @[PipelineReg.scala 23:25]
    .clock(imemrh_clock),
    .reset(imemrh_reset),
    .io_ren(imemrh_io_ren),
    .io_raddr(imemrh_io_raddr),
    .io_imem_raddr(imemrh_io_imem_raddr)
  );
  assign io_imem_addr = imemrh_io_imem_raddr; // @[PipelineReg.scala 27:21]
  assign io_pr_valid_out = valid; // @[PipelineReg.scala 29:21]
  assign io_pc_out = pc; // @[PipelineReg.scala 30:21]
  assign io_inst_out = io_imem_data; // @[PipelineReg.scala 31:21]
  assign imemrh_clock = clock;
  assign imemrh_reset = reset;
  assign imemrh_io_ren = io_pr_en; // @[PipelineReg.scala 24:21]
  assign imemrh_io_raddr = io_pc_in; // @[PipelineReg.scala 25:21]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 27:20]
      valid <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      valid <= io_pr_valid_in; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      pc <= 64'h7ffffffc; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      pc <= io_pc_in; // @[Reg.scala 28:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  pc = _RAND_1[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ExeReg(
  input         clock,
  input         reset,
  input         io_pr_valid_in,
  output        io_pr_valid_out,
  input         io_pr_en,
  input  [63:0] io_pc_in,
  input  [31:0] io_inst_in,
  input         io_rd_en_in,
  input  [4:0]  io_rd_addr_in,
  input  [63:0] io_imm_in,
  input  [63:0] io_op1_in,
  input  [63:0] io_op2_in,
  input  [4:0]  io_rs1_addr_in,
  input  [5:0]  io_decode_info_in_fu_code,
  input  [15:0] io_decode_info_in_alu_code,
  input  [7:0]  io_decode_info_in_bu_code,
  input  [6:0]  io_decode_info_in_lu_code,
  input  [3:0]  io_decode_info_in_su_code,
  input  [9:0]  io_decode_info_in_mdu_code,
  input  [6:0]  io_decode_info_in_csru_code,
  input         io_putch_in,
  output [63:0] io_pc_out,
  output [31:0] io_inst_out,
  output        io_rd_en_out,
  output [4:0]  io_rd_addr_out,
  output [63:0] io_imm_out,
  output [63:0] io_op1_out,
  output [63:0] io_op2_out,
  output [4:0]  io_rs1_addr_out,
  output [5:0]  io_decode_info_out_fu_code,
  output [15:0] io_decode_info_out_alu_code,
  output [7:0]  io_decode_info_out_bu_code,
  output [6:0]  io_decode_info_out_lu_code,
  output [3:0]  io_decode_info_out_su_code,
  output [9:0]  io_decode_info_out_mdu_code,
  output [6:0]  io_decode_info_out_csru_code,
  output        io_putch_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  reg  valid; // @[Reg.scala 27:20]
  reg [63:0] pc; // @[Reg.scala 27:20]
  reg [31:0] inst; // @[Reg.scala 27:20]
  reg  rd_en; // @[Reg.scala 27:20]
  reg [4:0] rd_addr; // @[Reg.scala 27:20]
  reg [63:0] imm; // @[Reg.scala 27:20]
  reg [63:0] op1; // @[Reg.scala 27:20]
  reg [63:0] op2; // @[Reg.scala 27:20]
  reg [5:0] fu_code; // @[Reg.scala 27:20]
  reg [15:0] alu_code; // @[Reg.scala 27:20]
  reg [7:0] bu_code; // @[Reg.scala 27:20]
  reg [6:0] lu_code; // @[Reg.scala 27:20]
  reg [3:0] su_code; // @[Reg.scala 27:20]
  reg [9:0] mdu_code; // @[Reg.scala 27:20]
  reg [6:0] csru_code; // @[Reg.scala 27:20]
  reg [4:0] io_rs1_addr_out_r; // @[Reg.scala 27:20]
  reg  io_putch_out_r; // @[Reg.scala 27:20]
  assign io_pr_valid_out = valid; // @[PipelineReg.scala 78:21]
  assign io_pc_out = pc; // @[PipelineReg.scala 79:15]
  assign io_inst_out = inst; // @[PipelineReg.scala 80:17]
  assign io_rd_en_out = rd_en; // @[PipelineReg.scala 81:18]
  assign io_rd_addr_out = rd_addr; // @[PipelineReg.scala 82:20]
  assign io_imm_out = imm; // @[PipelineReg.scala 83:16]
  assign io_op1_out = op1; // @[PipelineReg.scala 84:16]
  assign io_op2_out = op2; // @[PipelineReg.scala 85:16]
  assign io_rs1_addr_out = io_rs1_addr_out_r; // @[PipelineReg.scala 86:21]
  assign io_decode_info_out_fu_code = fu_code; // @[PipelineReg.scala 87:32]
  assign io_decode_info_out_alu_code = alu_code; // @[PipelineReg.scala 88:33]
  assign io_decode_info_out_bu_code = bu_code; // @[PipelineReg.scala 89:32]
  assign io_decode_info_out_lu_code = lu_code; // @[PipelineReg.scala 90:32]
  assign io_decode_info_out_su_code = su_code; // @[PipelineReg.scala 91:32]
  assign io_decode_info_out_mdu_code = mdu_code; // @[PipelineReg.scala 92:33]
  assign io_decode_info_out_csru_code = csru_code; // @[PipelineReg.scala 93:34]
  assign io_putch_out = io_putch_out_r; // @[PipelineReg.scala 95:18]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 27:20]
      valid <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      valid <= io_pr_valid_in; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      pc <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      pc <= io_pc_in; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      inst <= 32'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      inst <= io_inst_in; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      rd_en <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      rd_en <= io_rd_en_in; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      rd_addr <= 5'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      rd_addr <= io_rd_addr_in; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      imm <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      imm <= io_imm_in; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      op1 <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      op1 <= io_op1_in; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      op2 <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      op2 <= io_op2_in; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      fu_code <= 6'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      fu_code <= io_decode_info_in_fu_code; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      alu_code <= 16'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      alu_code <= io_decode_info_in_alu_code; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      bu_code <= 8'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      bu_code <= io_decode_info_in_bu_code; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      lu_code <= 7'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      lu_code <= io_decode_info_in_lu_code; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      su_code <= 4'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      su_code <= io_decode_info_in_su_code; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      mdu_code <= 10'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      mdu_code <= io_decode_info_in_mdu_code; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      csru_code <= 7'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      csru_code <= io_decode_info_in_csru_code; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      io_rs1_addr_out_r <= 5'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      io_rs1_addr_out_r <= io_rs1_addr_in; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      io_putch_out_r <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      io_putch_out_r <= io_putch_in; // @[Reg.scala 28:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  pc = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  inst = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  rd_en = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  rd_addr = _RAND_4[4:0];
  _RAND_5 = {2{`RANDOM}};
  imm = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  op1 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  op2 = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  fu_code = _RAND_8[5:0];
  _RAND_9 = {1{`RANDOM}};
  alu_code = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  bu_code = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  lu_code = _RAND_11[6:0];
  _RAND_12 = {1{`RANDOM}};
  su_code = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  mdu_code = _RAND_13[9:0];
  _RAND_14 = {1{`RANDOM}};
  csru_code = _RAND_14[6:0];
  _RAND_15 = {1{`RANDOM}};
  io_rs1_addr_out_r = _RAND_15[4:0];
  _RAND_16 = {1{`RANDOM}};
  io_putch_out_r = _RAND_16[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MemReg(
  input         clock,
  input         reset,
  input         io_pr_valid_in,
  output        io_pr_valid_out,
  input         io_pr_en,
  input  [63:0] io_pc_in,
  input  [31:0] io_inst_in,
  input         io_rd_en_in,
  input  [4:0]  io_rd_addr_in,
  input  [63:0] io_alu_out_in,
  input  [63:0] io_bu_out_in,
  input  [63:0] io_mdu_out_in,
  input  [63:0] io_csru_out_in,
  input  [63:0] io_imm_in,
  input  [63:0] io_op1_in,
  input  [63:0] io_op2_in,
  input  [5:0]  io_decode_info_in_fu_code,
  input  [6:0]  io_decode_info_in_lu_code,
  input  [3:0]  io_decode_info_in_su_code,
  input  [6:0]  io_decode_info_in_csru_code,
  input         io_putch_in,
  input         io_csr_wen_in,
  input  [11:0] io_csr_waddr_in,
  input  [63:0] io_csr_wdata_in,
  output [63:0] io_pc_out,
  output [31:0] io_inst_out,
  output        io_rd_en_out,
  output [4:0]  io_rd_addr_out,
  output [63:0] io_alu_out_out,
  output [63:0] io_bu_out_out,
  output [63:0] io_mdu_out_out,
  output [63:0] io_csru_out_out,
  output [63:0] io_imm_out,
  output [63:0] io_op1_out,
  output [63:0] io_op2_out,
  output [5:0]  io_decode_info_out_fu_code,
  output [6:0]  io_decode_info_out_lu_code,
  output [3:0]  io_decode_info_out_su_code,
  output [6:0]  io_decode_info_out_csru_code,
  output        io_putch_out,
  output        io_csr_wen_out,
  output [11:0] io_csr_waddr_out,
  output [63:0] io_csr_wdata_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [63:0] _RAND_19;
`endif // RANDOMIZE_REG_INIT
  reg  valid; // @[Reg.scala 27:20]
  reg [63:0] pc; // @[Reg.scala 27:20]
  reg [31:0] inst; // @[Reg.scala 27:20]
  reg  rd_en; // @[Reg.scala 27:20]
  reg [4:0] rd_addr; // @[Reg.scala 27:20]
  reg [63:0] alu_out; // @[Reg.scala 27:20]
  reg [63:0] bu_out; // @[Reg.scala 27:20]
  reg [63:0] mdu_out; // @[Reg.scala 27:20]
  reg [63:0] csru_out; // @[Reg.scala 27:20]
  reg [63:0] imm; // @[Reg.scala 27:20]
  reg [63:0] op1; // @[Reg.scala 27:20]
  reg [63:0] op2; // @[Reg.scala 27:20]
  reg [5:0] fu_code; // @[Reg.scala 27:20]
  reg [6:0] lu_code; // @[Reg.scala 27:20]
  reg [3:0] su_code; // @[Reg.scala 27:20]
  reg [6:0] csru_code; // @[Reg.scala 27:20]
  reg  io_putch_out_r; // @[Reg.scala 27:20]
  reg  io_csr_wen_out_r; // @[Reg.scala 27:20]
  reg [11:0] io_csr_waddr_out_r; // @[Reg.scala 27:20]
  reg [63:0] io_csr_wdata_out_r; // @[Reg.scala 27:20]
  assign io_pr_valid_out = valid; // @[PipelineReg.scala 161:21]
  assign io_pc_out = pc; // @[PipelineReg.scala 162:15]
  assign io_inst_out = inst; // @[PipelineReg.scala 163:17]
  assign io_rd_en_out = rd_en; // @[PipelineReg.scala 164:18]
  assign io_rd_addr_out = rd_addr; // @[PipelineReg.scala 165:20]
  assign io_alu_out_out = alu_out; // @[PipelineReg.scala 166:20]
  assign io_bu_out_out = bu_out; // @[PipelineReg.scala 167:19]
  assign io_mdu_out_out = mdu_out; // @[PipelineReg.scala 168:20]
  assign io_csru_out_out = csru_out; // @[PipelineReg.scala 169:21]
  assign io_imm_out = imm; // @[PipelineReg.scala 171:16]
  assign io_op1_out = op1; // @[PipelineReg.scala 172:16]
  assign io_op2_out = op2; // @[PipelineReg.scala 173:16]
  assign io_decode_info_out_fu_code = fu_code; // @[PipelineReg.scala 174:32]
  assign io_decode_info_out_lu_code = lu_code; // @[PipelineReg.scala 177:32]
  assign io_decode_info_out_su_code = su_code; // @[PipelineReg.scala 178:32]
  assign io_decode_info_out_csru_code = csru_code; // @[PipelineReg.scala 180:34]
  assign io_putch_out = io_putch_out_r; // @[PipelineReg.scala 182:22]
  assign io_csr_wen_out = io_csr_wen_out_r; // @[PipelineReg.scala 183:22]
  assign io_csr_waddr_out = io_csr_waddr_out_r; // @[PipelineReg.scala 184:22]
  assign io_csr_wdata_out = io_csr_wdata_out_r; // @[PipelineReg.scala 185:22]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 27:20]
      valid <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      valid <= io_pr_valid_in; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      pc <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      pc <= io_pc_in; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      inst <= 32'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      inst <= io_inst_in; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      rd_en <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      rd_en <= io_rd_en_in; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      rd_addr <= 5'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      rd_addr <= io_rd_addr_in; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      alu_out <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      alu_out <= io_alu_out_in; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      bu_out <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      bu_out <= io_bu_out_in; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      mdu_out <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      mdu_out <= io_mdu_out_in; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      csru_out <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      csru_out <= io_csru_out_in; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      imm <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      imm <= io_imm_in; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      op1 <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      op1 <= io_op1_in; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      op2 <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      op2 <= io_op2_in; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      fu_code <= 6'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      fu_code <= io_decode_info_in_fu_code; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      lu_code <= 7'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      lu_code <= io_decode_info_in_lu_code; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      su_code <= 4'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      su_code <= io_decode_info_in_su_code; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      csru_code <= 7'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      csru_code <= io_decode_info_in_csru_code; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      io_putch_out_r <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      io_putch_out_r <= io_putch_in; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      io_csr_wen_out_r <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      io_csr_wen_out_r <= io_csr_wen_in; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      io_csr_waddr_out_r <= 12'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      io_csr_waddr_out_r <= io_csr_waddr_in; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      io_csr_wdata_out_r <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      io_csr_wdata_out_r <= io_csr_wdata_in; // @[Reg.scala 28:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  pc = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  inst = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  rd_en = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  rd_addr = _RAND_4[4:0];
  _RAND_5 = {2{`RANDOM}};
  alu_out = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  bu_out = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  mdu_out = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  csru_out = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  imm = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  op1 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  op2 = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  fu_code = _RAND_12[5:0];
  _RAND_13 = {1{`RANDOM}};
  lu_code = _RAND_13[6:0];
  _RAND_14 = {1{`RANDOM}};
  su_code = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  csru_code = _RAND_15[6:0];
  _RAND_16 = {1{`RANDOM}};
  io_putch_out_r = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  io_csr_wen_out_r = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  io_csr_waddr_out_r = _RAND_18[11:0];
  _RAND_19 = {2{`RANDOM}};
  io_csr_wdata_out_r = _RAND_19[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module WBReg(
  input         clock,
  input         reset,
  input         io_pr_valid_in,
  output        io_pr_valid_out,
  input         io_pr_en,
  input  [63:0] io_pc_in,
  input  [31:0] io_inst_in,
  input         io_rd_en_in,
  input  [4:0]  io_rd_addr_in,
  input  [63:0] io_alu_out_in,
  input  [63:0] io_bu_out_in,
  input  [63:0] io_mdu_out_in,
  input  [63:0] io_csru_out_in,
  input  [5:0]  io_fu_code_in,
  input  [6:0]  io_lu_code_in,
  input  [6:0]  io_csru_code_in,
  input  [5:0]  io_lu_shift_in,
  input         io_putch_in,
  input         io_csr_wen_in,
  input  [11:0] io_csr_waddr_in,
  input  [63:0] io_csr_wdata_in,
  output [63:0] io_pc_out,
  output [31:0] io_inst_out,
  output        io_rd_en_out,
  output [4:0]  io_rd_addr_out,
  output [63:0] io_alu_out_out,
  output [63:0] io_bu_out_out,
  output [63:0] io_mdu_out_out,
  output [63:0] io_csru_out_out,
  output [5:0]  io_fu_code_out,
  output [6:0]  io_lu_code_out,
  output [6:0]  io_csru_code_out,
  output [5:0]  io_lu_shift_out,
  output        io_putch_out,
  output        io_csr_wen_out,
  output [11:0] io_csr_waddr_out,
  output [63:0] io_csr_wdata_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [63:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  reg  valid; // @[Reg.scala 27:20]
  reg [63:0] pc; // @[Reg.scala 27:20]
  reg [31:0] inst; // @[Reg.scala 27:20]
  reg  rd_en; // @[Reg.scala 27:20]
  reg [4:0] rd_addr; // @[Reg.scala 27:20]
  reg [63:0] alu_out; // @[Reg.scala 27:20]
  reg [63:0] bu_out; // @[Reg.scala 27:20]
  reg [63:0] mdu_out; // @[Reg.scala 27:20]
  reg [63:0] csru_out; // @[Reg.scala 27:20]
  reg [5:0] fu_code; // @[Reg.scala 27:20]
  reg [6:0] lu_code; // @[Reg.scala 27:20]
  reg [6:0] csru_code; // @[Reg.scala 27:20]
  reg [5:0] lu_shift; // @[Reg.scala 27:20]
  reg  io_putch_out_r; // @[Reg.scala 27:20]
  reg  io_csr_wen_out_r; // @[Reg.scala 27:20]
  reg [11:0] io_csr_waddr_out_r; // @[Reg.scala 27:20]
  reg [63:0] io_csr_wdata_out_r; // @[Reg.scala 27:20]
  assign io_pr_valid_out = valid; // @[PipelineReg.scala 246:21]
  assign io_pc_out = pc; // @[PipelineReg.scala 247:15]
  assign io_inst_out = inst; // @[PipelineReg.scala 248:17]
  assign io_rd_en_out = rd_en; // @[PipelineReg.scala 249:18]
  assign io_rd_addr_out = rd_addr; // @[PipelineReg.scala 250:20]
  assign io_alu_out_out = alu_out; // @[PipelineReg.scala 251:20]
  assign io_bu_out_out = bu_out; // @[PipelineReg.scala 252:19]
  assign io_mdu_out_out = mdu_out; // @[PipelineReg.scala 253:20]
  assign io_csru_out_out = csru_out; // @[PipelineReg.scala 254:21]
  assign io_fu_code_out = fu_code; // @[PipelineReg.scala 256:20]
  assign io_lu_code_out = lu_code; // @[PipelineReg.scala 257:20]
  assign io_csru_code_out = csru_code; // @[PipelineReg.scala 258:22]
  assign io_lu_shift_out = lu_shift; // @[PipelineReg.scala 259:21]
  assign io_putch_out = io_putch_out_r; // @[PipelineReg.scala 261:18]
  assign io_csr_wen_out = io_csr_wen_out_r; // @[PipelineReg.scala 262:22]
  assign io_csr_waddr_out = io_csr_waddr_out_r; // @[PipelineReg.scala 263:22]
  assign io_csr_wdata_out = io_csr_wdata_out_r; // @[PipelineReg.scala 264:22]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 27:20]
      valid <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      valid <= io_pr_valid_in; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      pc <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      pc <= io_pc_in; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      inst <= 32'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      inst <= io_inst_in; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      rd_en <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      rd_en <= io_rd_en_in; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      rd_addr <= 5'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      rd_addr <= io_rd_addr_in; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      alu_out <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      alu_out <= io_alu_out_in; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      bu_out <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      bu_out <= io_bu_out_in; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      mdu_out <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      mdu_out <= io_mdu_out_in; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      csru_out <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      csru_out <= io_csru_out_in; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      fu_code <= 6'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      fu_code <= io_fu_code_in; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      lu_code <= 7'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      lu_code <= io_lu_code_in; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      csru_code <= 7'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      csru_code <= io_csru_code_in; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      lu_shift <= 6'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      lu_shift <= io_lu_shift_in; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      io_putch_out_r <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      io_putch_out_r <= io_putch_in; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      io_csr_wen_out_r <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      io_csr_wen_out_r <= io_csr_wen_in; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      io_csr_waddr_out_r <= 12'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      io_csr_waddr_out_r <= io_csr_waddr_in; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      io_csr_wdata_out_r <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_pr_en) begin // @[Reg.scala 28:19]
      io_csr_wdata_out_r <= io_csr_wdata_in; // @[Reg.scala 28:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  pc = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  inst = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  rd_en = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  rd_addr = _RAND_4[4:0];
  _RAND_5 = {2{`RANDOM}};
  alu_out = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  bu_out = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  mdu_out = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  csru_out = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  fu_code = _RAND_9[5:0];
  _RAND_10 = {1{`RANDOM}};
  lu_code = _RAND_10[6:0];
  _RAND_11 = {1{`RANDOM}};
  csru_code = _RAND_11[6:0];
  _RAND_12 = {1{`RANDOM}};
  lu_shift = _RAND_12[5:0];
  _RAND_13 = {1{`RANDOM}};
  io_putch_out_r = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  io_csr_wen_out_r = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  io_csr_waddr_out_r = _RAND_15[11:0];
  _RAND_16 = {2{`RANDOM}};
  io_csr_wdata_out_r = _RAND_16[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Core(
  input         clock,
  input         reset,
  output [63:0] io_imem_addr,
  input  [31:0] io_imem_data,
  input         io_imem_data_ok,
  output        io_dmem_en,
  output        io_dmem_op,
  output [63:0] io_dmem_addr,
  output [63:0] io_dmem_wdata,
  output [7:0]  io_dmem_wmask,
  input         io_dmem_ok,
  input  [63:0] io_dmem_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire  ifu_reset; // @[Core.scala 28:23]
  wire  ifu_io_jump_en; // @[Core.scala 28:23]
  wire [63:0] ifu_io_jump_pc; // @[Core.scala 28:23]
  wire  ifu_io_en; // @[Core.scala 28:23]
  wire [63:0] ifu_io_pc; // @[Core.scala 28:23]
  wire [63:0] ifu_io_next_pc; // @[Core.scala 28:23]
  wire  ifu_io_valid; // @[Core.scala 28:23]
  wire [63:0] idu_io_pc; // @[Core.scala 29:23]
  wire [31:0] idu_io_inst; // @[Core.scala 29:23]
  wire  idu_io_rs1_en; // @[Core.scala 29:23]
  wire  idu_io_rs2_en; // @[Core.scala 29:23]
  wire [4:0] idu_io_rs1_addr; // @[Core.scala 29:23]
  wire [4:0] idu_io_rs2_addr; // @[Core.scala 29:23]
  wire [63:0] idu_io_rs1_data; // @[Core.scala 29:23]
  wire [63:0] idu_io_rs2_data; // @[Core.scala 29:23]
  wire  idu_io_rd_en; // @[Core.scala 29:23]
  wire [4:0] idu_io_rd_addr; // @[Core.scala 29:23]
  wire [5:0] idu_io_decode_info_fu_code; // @[Core.scala 29:23]
  wire [15:0] idu_io_decode_info_alu_code; // @[Core.scala 29:23]
  wire [7:0] idu_io_decode_info_bu_code; // @[Core.scala 29:23]
  wire [6:0] idu_io_decode_info_lu_code; // @[Core.scala 29:23]
  wire [3:0] idu_io_decode_info_su_code; // @[Core.scala 29:23]
  wire [9:0] idu_io_decode_info_mdu_code; // @[Core.scala 29:23]
  wire [6:0] idu_io_decode_info_csru_code; // @[Core.scala 29:23]
  wire  idu_io_jump_en; // @[Core.scala 29:23]
  wire [63:0] idu_io_jump_pc; // @[Core.scala 29:23]
  wire [63:0] idu_io_op1; // @[Core.scala 29:23]
  wire [63:0] idu_io_op2; // @[Core.scala 29:23]
  wire [63:0] idu_io_imm; // @[Core.scala 29:23]
  wire  idu_io_putch; // @[Core.scala 29:23]
  wire [63:0] idu_io_mtvec; // @[Core.scala 29:23]
  wire [63:0] idu_io_mepc; // @[Core.scala 29:23]
  wire [15:0] ieu_io_decode_info_alu_code; // @[Core.scala 30:23]
  wire [7:0] ieu_io_decode_info_bu_code; // @[Core.scala 30:23]
  wire [9:0] ieu_io_decode_info_mdu_code; // @[Core.scala 30:23]
  wire [6:0] ieu_io_decode_info_csru_code; // @[Core.scala 30:23]
  wire [63:0] ieu_io_op1; // @[Core.scala 30:23]
  wire [63:0] ieu_io_op2; // @[Core.scala 30:23]
  wire [63:0] ieu_io_pc; // @[Core.scala 30:23]
  wire [63:0] ieu_io_alu_out; // @[Core.scala 30:23]
  wire [63:0] ieu_io_bu_out; // @[Core.scala 30:23]
  wire [63:0] ieu_io_mdu_out; // @[Core.scala 30:23]
  wire [63:0] ieu_io_csru_out; // @[Core.scala 30:23]
  wire [4:0] ieu_io_rs1_addr; // @[Core.scala 30:23]
  wire [11:0] ieu_io_csr_raddr; // @[Core.scala 30:23]
  wire [63:0] ieu_io_csr_rdata; // @[Core.scala 30:23]
  wire  ieu_io_csr_wen; // @[Core.scala 30:23]
  wire [11:0] ieu_io_csr_waddr; // @[Core.scala 30:23]
  wire [63:0] ieu_io_csr_wdata; // @[Core.scala 30:23]
  wire  rfu_clock; // @[Core.scala 31:23]
  wire  rfu_reset; // @[Core.scala 31:23]
  wire [4:0] rfu_io_rs1_addr; // @[Core.scala 31:23]
  wire [4:0] rfu_io_rs2_addr; // @[Core.scala 31:23]
  wire [63:0] rfu_io_rs1_data; // @[Core.scala 31:23]
  wire [63:0] rfu_io_rs2_data; // @[Core.scala 31:23]
  wire [4:0] rfu_io_rd_addr; // @[Core.scala 31:23]
  wire [63:0] rfu_io_rd_data; // @[Core.scala 31:23]
  wire  rfu_io_rd_en; // @[Core.scala 31:23]
  wire [63:0] rfu_rf_10; // @[Core.scala 31:23]
  wire  csru_clock; // @[Core.scala 32:23]
  wire  csru_reset; // @[Core.scala 32:23]
  wire [11:0] csru_io_raddr; // @[Core.scala 32:23]
  wire [63:0] csru_io_rdata; // @[Core.scala 32:23]
  wire  csru_io_wen; // @[Core.scala 32:23]
  wire [11:0] csru_io_waddr; // @[Core.scala 32:23]
  wire [63:0] csru_io_wdata; // @[Core.scala 32:23]
  wire  csru_io_csru_code_valid; // @[Core.scala 32:23]
  wire [6:0] csru_io_csru_code; // @[Core.scala 32:23]
  wire [63:0] csru_io_pc; // @[Core.scala 32:23]
  wire [63:0] csru_io_mtvec; // @[Core.scala 32:23]
  wire [63:0] csru_io_mepc; // @[Core.scala 32:23]
  wire [6:0] preamu_io_lu_code; // @[Core.scala 33:23]
  wire [3:0] preamu_io_su_code; // @[Core.scala 33:23]
  wire [63:0] preamu_io_op1; // @[Core.scala 33:23]
  wire [63:0] preamu_io_op2; // @[Core.scala 33:23]
  wire [63:0] preamu_io_imm; // @[Core.scala 33:23]
  wire [5:0] preamu_io_lu_shift; // @[Core.scala 33:23]
  wire  preamu_io_ren; // @[Core.scala 33:23]
  wire [63:0] preamu_io_raddr; // @[Core.scala 33:23]
  wire  preamu_io_wen; // @[Core.scala 33:23]
  wire [63:0] preamu_io_waddr; // @[Core.scala 33:23]
  wire [63:0] preamu_io_wdata; // @[Core.scala 33:23]
  wire [7:0] preamu_io_wmask; // @[Core.scala 33:23]
  wire [6:0] amu_io_lu_code; // @[Core.scala 34:23]
  wire [5:0] amu_io_lu_shift; // @[Core.scala 34:23]
  wire [63:0] amu_io_rdata; // @[Core.scala 34:23]
  wire [63:0] amu_io_lu_out; // @[Core.scala 34:23]
  wire [5:0] wbu_io_fu_code; // @[Core.scala 35:23]
  wire [63:0] wbu_io_alu_out; // @[Core.scala 35:23]
  wire [63:0] wbu_io_bu_out; // @[Core.scala 35:23]
  wire [63:0] wbu_io_mdu_out; // @[Core.scala 35:23]
  wire [63:0] wbu_io_lu_out; // @[Core.scala 35:23]
  wire [63:0] wbu_io_csru_out; // @[Core.scala 35:23]
  wire [63:0] wbu_io_out; // @[Core.scala 35:23]
  wire  rfconflict_io_rs_valid; // @[Core.scala 37:27]
  wire  rfconflict_io_rs1_en; // @[Core.scala 37:27]
  wire  rfconflict_io_rs2_en; // @[Core.scala 37:27]
  wire [4:0] rfconflict_io_rs1_addr; // @[Core.scala 37:27]
  wire [4:0] rfconflict_io_rs2_addr; // @[Core.scala 37:27]
  wire  rfconflict_io_rd1_valid; // @[Core.scala 37:27]
  wire  rfconflict_io_rd1_en; // @[Core.scala 37:27]
  wire [4:0] rfconflict_io_rd1_addr; // @[Core.scala 37:27]
  wire  rfconflict_io_rd2_valid; // @[Core.scala 37:27]
  wire  rfconflict_io_rd2_en; // @[Core.scala 37:27]
  wire [4:0] rfconflict_io_rd2_addr; // @[Core.scala 37:27]
  wire  rfconflict_io_rd3_valid; // @[Core.scala 37:27]
  wire  rfconflict_io_rd3_en; // @[Core.scala 37:27]
  wire [4:0] rfconflict_io_rd3_addr; // @[Core.scala 37:27]
  wire  rfconflict_io_conflict; // @[Core.scala 37:27]
  wire  idreg_clock; // @[Core.scala 39:23]
  wire  idreg_reset; // @[Core.scala 39:23]
  wire [63:0] idreg_io_imem_addr; // @[Core.scala 39:23]
  wire [31:0] idreg_io_imem_data; // @[Core.scala 39:23]
  wire  idreg_io_pr_valid_in; // @[Core.scala 39:23]
  wire  idreg_io_pr_valid_out; // @[Core.scala 39:23]
  wire  idreg_io_pr_en; // @[Core.scala 39:23]
  wire [63:0] idreg_io_pc_in; // @[Core.scala 39:23]
  wire [63:0] idreg_io_pc_out; // @[Core.scala 39:23]
  wire [31:0] idreg_io_inst_out; // @[Core.scala 39:23]
  wire  exereg_clock; // @[Core.scala 40:23]
  wire  exereg_reset; // @[Core.scala 40:23]
  wire  exereg_io_pr_valid_in; // @[Core.scala 40:23]
  wire  exereg_io_pr_valid_out; // @[Core.scala 40:23]
  wire  exereg_io_pr_en; // @[Core.scala 40:23]
  wire [63:0] exereg_io_pc_in; // @[Core.scala 40:23]
  wire [31:0] exereg_io_inst_in; // @[Core.scala 40:23]
  wire  exereg_io_rd_en_in; // @[Core.scala 40:23]
  wire [4:0] exereg_io_rd_addr_in; // @[Core.scala 40:23]
  wire [63:0] exereg_io_imm_in; // @[Core.scala 40:23]
  wire [63:0] exereg_io_op1_in; // @[Core.scala 40:23]
  wire [63:0] exereg_io_op2_in; // @[Core.scala 40:23]
  wire [4:0] exereg_io_rs1_addr_in; // @[Core.scala 40:23]
  wire [5:0] exereg_io_decode_info_in_fu_code; // @[Core.scala 40:23]
  wire [15:0] exereg_io_decode_info_in_alu_code; // @[Core.scala 40:23]
  wire [7:0] exereg_io_decode_info_in_bu_code; // @[Core.scala 40:23]
  wire [6:0] exereg_io_decode_info_in_lu_code; // @[Core.scala 40:23]
  wire [3:0] exereg_io_decode_info_in_su_code; // @[Core.scala 40:23]
  wire [9:0] exereg_io_decode_info_in_mdu_code; // @[Core.scala 40:23]
  wire [6:0] exereg_io_decode_info_in_csru_code; // @[Core.scala 40:23]
  wire  exereg_io_putch_in; // @[Core.scala 40:23]
  wire [63:0] exereg_io_pc_out; // @[Core.scala 40:23]
  wire [31:0] exereg_io_inst_out; // @[Core.scala 40:23]
  wire  exereg_io_rd_en_out; // @[Core.scala 40:23]
  wire [4:0] exereg_io_rd_addr_out; // @[Core.scala 40:23]
  wire [63:0] exereg_io_imm_out; // @[Core.scala 40:23]
  wire [63:0] exereg_io_op1_out; // @[Core.scala 40:23]
  wire [63:0] exereg_io_op2_out; // @[Core.scala 40:23]
  wire [4:0] exereg_io_rs1_addr_out; // @[Core.scala 40:23]
  wire [5:0] exereg_io_decode_info_out_fu_code; // @[Core.scala 40:23]
  wire [15:0] exereg_io_decode_info_out_alu_code; // @[Core.scala 40:23]
  wire [7:0] exereg_io_decode_info_out_bu_code; // @[Core.scala 40:23]
  wire [6:0] exereg_io_decode_info_out_lu_code; // @[Core.scala 40:23]
  wire [3:0] exereg_io_decode_info_out_su_code; // @[Core.scala 40:23]
  wire [9:0] exereg_io_decode_info_out_mdu_code; // @[Core.scala 40:23]
  wire [6:0] exereg_io_decode_info_out_csru_code; // @[Core.scala 40:23]
  wire  exereg_io_putch_out; // @[Core.scala 40:23]
  wire  memreg_clock; // @[Core.scala 41:23]
  wire  memreg_reset; // @[Core.scala 41:23]
  wire  memreg_io_pr_valid_in; // @[Core.scala 41:23]
  wire  memreg_io_pr_valid_out; // @[Core.scala 41:23]
  wire  memreg_io_pr_en; // @[Core.scala 41:23]
  wire [63:0] memreg_io_pc_in; // @[Core.scala 41:23]
  wire [31:0] memreg_io_inst_in; // @[Core.scala 41:23]
  wire  memreg_io_rd_en_in; // @[Core.scala 41:23]
  wire [4:0] memreg_io_rd_addr_in; // @[Core.scala 41:23]
  wire [63:0] memreg_io_alu_out_in; // @[Core.scala 41:23]
  wire [63:0] memreg_io_bu_out_in; // @[Core.scala 41:23]
  wire [63:0] memreg_io_mdu_out_in; // @[Core.scala 41:23]
  wire [63:0] memreg_io_csru_out_in; // @[Core.scala 41:23]
  wire [63:0] memreg_io_imm_in; // @[Core.scala 41:23]
  wire [63:0] memreg_io_op1_in; // @[Core.scala 41:23]
  wire [63:0] memreg_io_op2_in; // @[Core.scala 41:23]
  wire [5:0] memreg_io_decode_info_in_fu_code; // @[Core.scala 41:23]
  wire [6:0] memreg_io_decode_info_in_lu_code; // @[Core.scala 41:23]
  wire [3:0] memreg_io_decode_info_in_su_code; // @[Core.scala 41:23]
  wire [6:0] memreg_io_decode_info_in_csru_code; // @[Core.scala 41:23]
  wire  memreg_io_putch_in; // @[Core.scala 41:23]
  wire  memreg_io_csr_wen_in; // @[Core.scala 41:23]
  wire [11:0] memreg_io_csr_waddr_in; // @[Core.scala 41:23]
  wire [63:0] memreg_io_csr_wdata_in; // @[Core.scala 41:23]
  wire [63:0] memreg_io_pc_out; // @[Core.scala 41:23]
  wire [31:0] memreg_io_inst_out; // @[Core.scala 41:23]
  wire  memreg_io_rd_en_out; // @[Core.scala 41:23]
  wire [4:0] memreg_io_rd_addr_out; // @[Core.scala 41:23]
  wire [63:0] memreg_io_alu_out_out; // @[Core.scala 41:23]
  wire [63:0] memreg_io_bu_out_out; // @[Core.scala 41:23]
  wire [63:0] memreg_io_mdu_out_out; // @[Core.scala 41:23]
  wire [63:0] memreg_io_csru_out_out; // @[Core.scala 41:23]
  wire [63:0] memreg_io_imm_out; // @[Core.scala 41:23]
  wire [63:0] memreg_io_op1_out; // @[Core.scala 41:23]
  wire [63:0] memreg_io_op2_out; // @[Core.scala 41:23]
  wire [5:0] memreg_io_decode_info_out_fu_code; // @[Core.scala 41:23]
  wire [6:0] memreg_io_decode_info_out_lu_code; // @[Core.scala 41:23]
  wire [3:0] memreg_io_decode_info_out_su_code; // @[Core.scala 41:23]
  wire [6:0] memreg_io_decode_info_out_csru_code; // @[Core.scala 41:23]
  wire  memreg_io_putch_out; // @[Core.scala 41:23]
  wire  memreg_io_csr_wen_out; // @[Core.scala 41:23]
  wire [11:0] memreg_io_csr_waddr_out; // @[Core.scala 41:23]
  wire [63:0] memreg_io_csr_wdata_out; // @[Core.scala 41:23]
  wire  wbreg_clock; // @[Core.scala 42:23]
  wire  wbreg_reset; // @[Core.scala 42:23]
  wire  wbreg_io_pr_valid_in; // @[Core.scala 42:23]
  wire  wbreg_io_pr_valid_out; // @[Core.scala 42:23]
  wire  wbreg_io_pr_en; // @[Core.scala 42:23]
  wire [63:0] wbreg_io_pc_in; // @[Core.scala 42:23]
  wire [31:0] wbreg_io_inst_in; // @[Core.scala 42:23]
  wire  wbreg_io_rd_en_in; // @[Core.scala 42:23]
  wire [4:0] wbreg_io_rd_addr_in; // @[Core.scala 42:23]
  wire [63:0] wbreg_io_alu_out_in; // @[Core.scala 42:23]
  wire [63:0] wbreg_io_bu_out_in; // @[Core.scala 42:23]
  wire [63:0] wbreg_io_mdu_out_in; // @[Core.scala 42:23]
  wire [63:0] wbreg_io_csru_out_in; // @[Core.scala 42:23]
  wire [5:0] wbreg_io_fu_code_in; // @[Core.scala 42:23]
  wire [6:0] wbreg_io_lu_code_in; // @[Core.scala 42:23]
  wire [6:0] wbreg_io_csru_code_in; // @[Core.scala 42:23]
  wire [5:0] wbreg_io_lu_shift_in; // @[Core.scala 42:23]
  wire  wbreg_io_putch_in; // @[Core.scala 42:23]
  wire  wbreg_io_csr_wen_in; // @[Core.scala 42:23]
  wire [11:0] wbreg_io_csr_waddr_in; // @[Core.scala 42:23]
  wire [63:0] wbreg_io_csr_wdata_in; // @[Core.scala 42:23]
  wire [63:0] wbreg_io_pc_out; // @[Core.scala 42:23]
  wire [31:0] wbreg_io_inst_out; // @[Core.scala 42:23]
  wire  wbreg_io_rd_en_out; // @[Core.scala 42:23]
  wire [4:0] wbreg_io_rd_addr_out; // @[Core.scala 42:23]
  wire [63:0] wbreg_io_alu_out_out; // @[Core.scala 42:23]
  wire [63:0] wbreg_io_bu_out_out; // @[Core.scala 42:23]
  wire [63:0] wbreg_io_mdu_out_out; // @[Core.scala 42:23]
  wire [63:0] wbreg_io_csru_out_out; // @[Core.scala 42:23]
  wire [5:0] wbreg_io_fu_code_out; // @[Core.scala 42:23]
  wire [6:0] wbreg_io_lu_code_out; // @[Core.scala 42:23]
  wire [6:0] wbreg_io_csru_code_out; // @[Core.scala 42:23]
  wire [5:0] wbreg_io_lu_shift_out; // @[Core.scala 42:23]
  wire  wbreg_io_putch_out; // @[Core.scala 42:23]
  wire  wbreg_io_csr_wen_out; // @[Core.scala 42:23]
  wire [11:0] wbreg_io_csr_waddr_out; // @[Core.scala 42:23]
  wire [63:0] wbreg_io_csr_wdata_out; // @[Core.scala 42:23]
  wire  dt_ic_clock; // @[Core.scala 224:21]
  wire [7:0] dt_ic_coreid; // @[Core.scala 224:21]
  wire [7:0] dt_ic_index; // @[Core.scala 224:21]
  wire  dt_ic_valid; // @[Core.scala 224:21]
  wire [63:0] dt_ic_pc; // @[Core.scala 224:21]
  wire [31:0] dt_ic_instr; // @[Core.scala 224:21]
  wire [7:0] dt_ic_special; // @[Core.scala 224:21]
  wire  dt_ic_skip; // @[Core.scala 224:21]
  wire  dt_ic_isRVC; // @[Core.scala 224:21]
  wire  dt_ic_scFailed; // @[Core.scala 224:21]
  wire  dt_ic_wen; // @[Core.scala 224:21]
  wire [63:0] dt_ic_wdata; // @[Core.scala 224:21]
  wire [7:0] dt_ic_wdest; // @[Core.scala 224:21]
  wire  dt_ae_clock; // @[Core.scala 239:21]
  wire [7:0] dt_ae_coreid; // @[Core.scala 239:21]
  wire [31:0] dt_ae_intrNO; // @[Core.scala 239:21]
  wire [31:0] dt_ae_cause; // @[Core.scala 239:21]
  wire [63:0] dt_ae_exceptionPC; // @[Core.scala 239:21]
  wire [31:0] dt_ae_exceptionInst; // @[Core.scala 239:21]
  wire  dt_te_clock; // @[Core.scala 255:21]
  wire [7:0] dt_te_coreid; // @[Core.scala 255:21]
  wire  dt_te_valid; // @[Core.scala 255:21]
  wire [2:0] dt_te_code; // @[Core.scala 255:21]
  wire [63:0] dt_te_pc; // @[Core.scala 255:21]
  wire [63:0] dt_te_cycleCnt; // @[Core.scala 255:21]
  wire [63:0] dt_te_instrCnt; // @[Core.scala 255:21]
  wire  dmem_en = preamu_io_ren | preamu_io_wen; // @[Core.scala 106:31]
  wire  imem_not_ok = ~io_imem_data_ok; // @[Core.scala 178:21]
  wire  dmem_not_ok = ~io_dmem_ok; // @[Core.scala 179:21]
  wire  stall = rfconflict_io_conflict | imem_not_ok; // @[Core.scala 181:38]
  wire  _exereg_io_pr_valid_in_T = ~stall; // @[Core.scala 193:54]
  wire  _commit_valid_T = ~dmem_not_ok; // @[Core.scala 196:47]
  wire  commit_valid = wbreg_io_pr_valid_out & ~dmem_not_ok; // @[Core.scala 196:44]
  wire [31:0] _read_mcycle_T = wbreg_io_inst_out & 32'hfff0307f; // @[Core.scala 219:27]
  wire  read_mcycle = _read_mcycle_T == 32'hb0002073; // @[Core.scala 219:44]
  wire  read_mtime = wbreg_io_inst_out == 32'hff86b683; // @[Core.scala 220:25]
  wire  write_mtimecmp = wbreg_io_inst_out == 32'hd7b023; // @[Core.scala 221:29]
  reg  dt_ic_io_valid_REG; // @[Core.scala 228:31]
  reg [63:0] dt_ic_io_pc_REG; // @[Core.scala 229:31]
  reg [31:0] dt_ic_io_instr_REG; // @[Core.scala 230:31]
  reg  dt_ic_io_skip_REG; // @[Core.scala 232:31]
  reg  dt_ic_io_wen_REG; // @[Core.scala 235:31]
  reg [63:0] dt_ic_io_wdata_REG; // @[Core.scala 236:31]
  reg [4:0] dt_ic_io_wdest_REG; // @[Core.scala 237:31]
  reg [63:0] cycle_cnt; // @[Core.scala 246:26]
  reg [63:0] instr_cnt; // @[Core.scala 247:26]
  wire [63:0] _cycle_cnt_T_1 = cycle_cnt + 64'h1; // @[Core.scala 249:26]
  wire [63:0] _instr_cnt_T_1 = instr_cnt + 64'h1; // @[Core.scala 250:44]
  wire [63:0] rf_a0_0 = rfu_rf_10;
  IFetch ifu ( // @[Core.scala 28:23]
    .reset(ifu_reset),
    .io_jump_en(ifu_io_jump_en),
    .io_jump_pc(ifu_io_jump_pc),
    .io_en(ifu_io_en),
    .io_pc(ifu_io_pc),
    .io_next_pc(ifu_io_next_pc),
    .io_valid(ifu_io_valid)
  );
  Decode idu ( // @[Core.scala 29:23]
    .io_pc(idu_io_pc),
    .io_inst(idu_io_inst),
    .io_rs1_en(idu_io_rs1_en),
    .io_rs2_en(idu_io_rs2_en),
    .io_rs1_addr(idu_io_rs1_addr),
    .io_rs2_addr(idu_io_rs2_addr),
    .io_rs1_data(idu_io_rs1_data),
    .io_rs2_data(idu_io_rs2_data),
    .io_rd_en(idu_io_rd_en),
    .io_rd_addr(idu_io_rd_addr),
    .io_decode_info_fu_code(idu_io_decode_info_fu_code),
    .io_decode_info_alu_code(idu_io_decode_info_alu_code),
    .io_decode_info_bu_code(idu_io_decode_info_bu_code),
    .io_decode_info_lu_code(idu_io_decode_info_lu_code),
    .io_decode_info_su_code(idu_io_decode_info_su_code),
    .io_decode_info_mdu_code(idu_io_decode_info_mdu_code),
    .io_decode_info_csru_code(idu_io_decode_info_csru_code),
    .io_jump_en(idu_io_jump_en),
    .io_jump_pc(idu_io_jump_pc),
    .io_op1(idu_io_op1),
    .io_op2(idu_io_op2),
    .io_imm(idu_io_imm),
    .io_putch(idu_io_putch),
    .io_mtvec(idu_io_mtvec),
    .io_mepc(idu_io_mepc)
  );
  Execution ieu ( // @[Core.scala 30:23]
    .io_decode_info_alu_code(ieu_io_decode_info_alu_code),
    .io_decode_info_bu_code(ieu_io_decode_info_bu_code),
    .io_decode_info_mdu_code(ieu_io_decode_info_mdu_code),
    .io_decode_info_csru_code(ieu_io_decode_info_csru_code),
    .io_op1(ieu_io_op1),
    .io_op2(ieu_io_op2),
    .io_pc(ieu_io_pc),
    .io_alu_out(ieu_io_alu_out),
    .io_bu_out(ieu_io_bu_out),
    .io_mdu_out(ieu_io_mdu_out),
    .io_csru_out(ieu_io_csru_out),
    .io_rs1_addr(ieu_io_rs1_addr),
    .io_csr_raddr(ieu_io_csr_raddr),
    .io_csr_rdata(ieu_io_csr_rdata),
    .io_csr_wen(ieu_io_csr_wen),
    .io_csr_waddr(ieu_io_csr_waddr),
    .io_csr_wdata(ieu_io_csr_wdata)
  );
  RegFile rfu ( // @[Core.scala 31:23]
    .clock(rfu_clock),
    .reset(rfu_reset),
    .io_rs1_addr(rfu_io_rs1_addr),
    .io_rs2_addr(rfu_io_rs2_addr),
    .io_rs1_data(rfu_io_rs1_data),
    .io_rs2_data(rfu_io_rs2_data),
    .io_rd_addr(rfu_io_rd_addr),
    .io_rd_data(rfu_io_rd_data),
    .io_rd_en(rfu_io_rd_en),
    .rf_10(rfu_rf_10)
  );
  Csr csru ( // @[Core.scala 32:23]
    .clock(csru_clock),
    .reset(csru_reset),
    .io_raddr(csru_io_raddr),
    .io_rdata(csru_io_rdata),
    .io_wen(csru_io_wen),
    .io_waddr(csru_io_waddr),
    .io_wdata(csru_io_wdata),
    .io_csru_code_valid(csru_io_csru_code_valid),
    .io_csru_code(csru_io_csru_code),
    .io_pc(csru_io_pc),
    .io_mtvec(csru_io_mtvec),
    .io_mepc(csru_io_mepc)
  );
  PreAccessMemory preamu ( // @[Core.scala 33:23]
    .io_lu_code(preamu_io_lu_code),
    .io_su_code(preamu_io_su_code),
    .io_op1(preamu_io_op1),
    .io_op2(preamu_io_op2),
    .io_imm(preamu_io_imm),
    .io_lu_shift(preamu_io_lu_shift),
    .io_ren(preamu_io_ren),
    .io_raddr(preamu_io_raddr),
    .io_wen(preamu_io_wen),
    .io_waddr(preamu_io_waddr),
    .io_wdata(preamu_io_wdata),
    .io_wmask(preamu_io_wmask)
  );
  AccessMemory amu ( // @[Core.scala 34:23]
    .io_lu_code(amu_io_lu_code),
    .io_lu_shift(amu_io_lu_shift),
    .io_rdata(amu_io_rdata),
    .io_lu_out(amu_io_lu_out)
  );
  WriteBack wbu ( // @[Core.scala 35:23]
    .io_fu_code(wbu_io_fu_code),
    .io_alu_out(wbu_io_alu_out),
    .io_bu_out(wbu_io_bu_out),
    .io_mdu_out(wbu_io_mdu_out),
    .io_lu_out(wbu_io_lu_out),
    .io_csru_out(wbu_io_csru_out),
    .io_out(wbu_io_out)
  );
  RegfileConflict rfconflict ( // @[Core.scala 37:27]
    .io_rs_valid(rfconflict_io_rs_valid),
    .io_rs1_en(rfconflict_io_rs1_en),
    .io_rs2_en(rfconflict_io_rs2_en),
    .io_rs1_addr(rfconflict_io_rs1_addr),
    .io_rs2_addr(rfconflict_io_rs2_addr),
    .io_rd1_valid(rfconflict_io_rd1_valid),
    .io_rd1_en(rfconflict_io_rd1_en),
    .io_rd1_addr(rfconflict_io_rd1_addr),
    .io_rd2_valid(rfconflict_io_rd2_valid),
    .io_rd2_en(rfconflict_io_rd2_en),
    .io_rd2_addr(rfconflict_io_rd2_addr),
    .io_rd3_valid(rfconflict_io_rd3_valid),
    .io_rd3_en(rfconflict_io_rd3_en),
    .io_rd3_addr(rfconflict_io_rd3_addr),
    .io_conflict(rfconflict_io_conflict)
  );
  IDReg idreg ( // @[Core.scala 39:23]
    .clock(idreg_clock),
    .reset(idreg_reset),
    .io_imem_addr(idreg_io_imem_addr),
    .io_imem_data(idreg_io_imem_data),
    .io_pr_valid_in(idreg_io_pr_valid_in),
    .io_pr_valid_out(idreg_io_pr_valid_out),
    .io_pr_en(idreg_io_pr_en),
    .io_pc_in(idreg_io_pc_in),
    .io_pc_out(idreg_io_pc_out),
    .io_inst_out(idreg_io_inst_out)
  );
  ExeReg exereg ( // @[Core.scala 40:23]
    .clock(exereg_clock),
    .reset(exereg_reset),
    .io_pr_valid_in(exereg_io_pr_valid_in),
    .io_pr_valid_out(exereg_io_pr_valid_out),
    .io_pr_en(exereg_io_pr_en),
    .io_pc_in(exereg_io_pc_in),
    .io_inst_in(exereg_io_inst_in),
    .io_rd_en_in(exereg_io_rd_en_in),
    .io_rd_addr_in(exereg_io_rd_addr_in),
    .io_imm_in(exereg_io_imm_in),
    .io_op1_in(exereg_io_op1_in),
    .io_op2_in(exereg_io_op2_in),
    .io_rs1_addr_in(exereg_io_rs1_addr_in),
    .io_decode_info_in_fu_code(exereg_io_decode_info_in_fu_code),
    .io_decode_info_in_alu_code(exereg_io_decode_info_in_alu_code),
    .io_decode_info_in_bu_code(exereg_io_decode_info_in_bu_code),
    .io_decode_info_in_lu_code(exereg_io_decode_info_in_lu_code),
    .io_decode_info_in_su_code(exereg_io_decode_info_in_su_code),
    .io_decode_info_in_mdu_code(exereg_io_decode_info_in_mdu_code),
    .io_decode_info_in_csru_code(exereg_io_decode_info_in_csru_code),
    .io_putch_in(exereg_io_putch_in),
    .io_pc_out(exereg_io_pc_out),
    .io_inst_out(exereg_io_inst_out),
    .io_rd_en_out(exereg_io_rd_en_out),
    .io_rd_addr_out(exereg_io_rd_addr_out),
    .io_imm_out(exereg_io_imm_out),
    .io_op1_out(exereg_io_op1_out),
    .io_op2_out(exereg_io_op2_out),
    .io_rs1_addr_out(exereg_io_rs1_addr_out),
    .io_decode_info_out_fu_code(exereg_io_decode_info_out_fu_code),
    .io_decode_info_out_alu_code(exereg_io_decode_info_out_alu_code),
    .io_decode_info_out_bu_code(exereg_io_decode_info_out_bu_code),
    .io_decode_info_out_lu_code(exereg_io_decode_info_out_lu_code),
    .io_decode_info_out_su_code(exereg_io_decode_info_out_su_code),
    .io_decode_info_out_mdu_code(exereg_io_decode_info_out_mdu_code),
    .io_decode_info_out_csru_code(exereg_io_decode_info_out_csru_code),
    .io_putch_out(exereg_io_putch_out)
  );
  MemReg memreg ( // @[Core.scala 41:23]
    .clock(memreg_clock),
    .reset(memreg_reset),
    .io_pr_valid_in(memreg_io_pr_valid_in),
    .io_pr_valid_out(memreg_io_pr_valid_out),
    .io_pr_en(memreg_io_pr_en),
    .io_pc_in(memreg_io_pc_in),
    .io_inst_in(memreg_io_inst_in),
    .io_rd_en_in(memreg_io_rd_en_in),
    .io_rd_addr_in(memreg_io_rd_addr_in),
    .io_alu_out_in(memreg_io_alu_out_in),
    .io_bu_out_in(memreg_io_bu_out_in),
    .io_mdu_out_in(memreg_io_mdu_out_in),
    .io_csru_out_in(memreg_io_csru_out_in),
    .io_imm_in(memreg_io_imm_in),
    .io_op1_in(memreg_io_op1_in),
    .io_op2_in(memreg_io_op2_in),
    .io_decode_info_in_fu_code(memreg_io_decode_info_in_fu_code),
    .io_decode_info_in_lu_code(memreg_io_decode_info_in_lu_code),
    .io_decode_info_in_su_code(memreg_io_decode_info_in_su_code),
    .io_decode_info_in_csru_code(memreg_io_decode_info_in_csru_code),
    .io_putch_in(memreg_io_putch_in),
    .io_csr_wen_in(memreg_io_csr_wen_in),
    .io_csr_waddr_in(memreg_io_csr_waddr_in),
    .io_csr_wdata_in(memreg_io_csr_wdata_in),
    .io_pc_out(memreg_io_pc_out),
    .io_inst_out(memreg_io_inst_out),
    .io_rd_en_out(memreg_io_rd_en_out),
    .io_rd_addr_out(memreg_io_rd_addr_out),
    .io_alu_out_out(memreg_io_alu_out_out),
    .io_bu_out_out(memreg_io_bu_out_out),
    .io_mdu_out_out(memreg_io_mdu_out_out),
    .io_csru_out_out(memreg_io_csru_out_out),
    .io_imm_out(memreg_io_imm_out),
    .io_op1_out(memreg_io_op1_out),
    .io_op2_out(memreg_io_op2_out),
    .io_decode_info_out_fu_code(memreg_io_decode_info_out_fu_code),
    .io_decode_info_out_lu_code(memreg_io_decode_info_out_lu_code),
    .io_decode_info_out_su_code(memreg_io_decode_info_out_su_code),
    .io_decode_info_out_csru_code(memreg_io_decode_info_out_csru_code),
    .io_putch_out(memreg_io_putch_out),
    .io_csr_wen_out(memreg_io_csr_wen_out),
    .io_csr_waddr_out(memreg_io_csr_waddr_out),
    .io_csr_wdata_out(memreg_io_csr_wdata_out)
  );
  WBReg wbreg ( // @[Core.scala 42:23]
    .clock(wbreg_clock),
    .reset(wbreg_reset),
    .io_pr_valid_in(wbreg_io_pr_valid_in),
    .io_pr_valid_out(wbreg_io_pr_valid_out),
    .io_pr_en(wbreg_io_pr_en),
    .io_pc_in(wbreg_io_pc_in),
    .io_inst_in(wbreg_io_inst_in),
    .io_rd_en_in(wbreg_io_rd_en_in),
    .io_rd_addr_in(wbreg_io_rd_addr_in),
    .io_alu_out_in(wbreg_io_alu_out_in),
    .io_bu_out_in(wbreg_io_bu_out_in),
    .io_mdu_out_in(wbreg_io_mdu_out_in),
    .io_csru_out_in(wbreg_io_csru_out_in),
    .io_fu_code_in(wbreg_io_fu_code_in),
    .io_lu_code_in(wbreg_io_lu_code_in),
    .io_csru_code_in(wbreg_io_csru_code_in),
    .io_lu_shift_in(wbreg_io_lu_shift_in),
    .io_putch_in(wbreg_io_putch_in),
    .io_csr_wen_in(wbreg_io_csr_wen_in),
    .io_csr_waddr_in(wbreg_io_csr_waddr_in),
    .io_csr_wdata_in(wbreg_io_csr_wdata_in),
    .io_pc_out(wbreg_io_pc_out),
    .io_inst_out(wbreg_io_inst_out),
    .io_rd_en_out(wbreg_io_rd_en_out),
    .io_rd_addr_out(wbreg_io_rd_addr_out),
    .io_alu_out_out(wbreg_io_alu_out_out),
    .io_bu_out_out(wbreg_io_bu_out_out),
    .io_mdu_out_out(wbreg_io_mdu_out_out),
    .io_csru_out_out(wbreg_io_csru_out_out),
    .io_fu_code_out(wbreg_io_fu_code_out),
    .io_lu_code_out(wbreg_io_lu_code_out),
    .io_csru_code_out(wbreg_io_csru_code_out),
    .io_lu_shift_out(wbreg_io_lu_shift_out),
    .io_putch_out(wbreg_io_putch_out),
    .io_csr_wen_out(wbreg_io_csr_wen_out),
    .io_csr_waddr_out(wbreg_io_csr_waddr_out),
    .io_csr_wdata_out(wbreg_io_csr_wdata_out)
  );
  DifftestInstrCommit dt_ic ( // @[Core.scala 224:21]
    .clock(dt_ic_clock),
    .coreid(dt_ic_coreid),
    .index(dt_ic_index),
    .valid(dt_ic_valid),
    .pc(dt_ic_pc),
    .instr(dt_ic_instr),
    .special(dt_ic_special),
    .skip(dt_ic_skip),
    .isRVC(dt_ic_isRVC),
    .scFailed(dt_ic_scFailed),
    .wen(dt_ic_wen),
    .wdata(dt_ic_wdata),
    .wdest(dt_ic_wdest)
  );
  DifftestArchEvent dt_ae ( // @[Core.scala 239:21]
    .clock(dt_ae_clock),
    .coreid(dt_ae_coreid),
    .intrNO(dt_ae_intrNO),
    .cause(dt_ae_cause),
    .exceptionPC(dt_ae_exceptionPC),
    .exceptionInst(dt_ae_exceptionInst)
  );
  DifftestTrapEvent dt_te ( // @[Core.scala 255:21]
    .clock(dt_te_clock),
    .coreid(dt_te_coreid),
    .valid(dt_te_valid),
    .code(dt_te_code),
    .pc(dt_te_pc),
    .cycleCnt(dt_te_cycleCnt),
    .instrCnt(dt_te_instrCnt)
  );
  assign io_imem_addr = idreg_io_imem_addr; // @[Core.scala 49:23]
  assign io_dmem_en = dmem_en & memreg_io_pr_valid_out; // @[Core.scala 109:28]
  assign io_dmem_op = preamu_io_wen; // @[Core.scala 110:17]
  assign io_dmem_addr = preamu_io_wen ? preamu_io_waddr : preamu_io_raddr; // @[Core.scala 108:22]
  assign io_dmem_wdata = preamu_io_wdata; // @[Core.scala 112:17]
  assign io_dmem_wmask = preamu_io_wmask; // @[Core.scala 113:17]
  assign ifu_reset = reset;
  assign ifu_io_jump_en = idu_io_jump_en; // @[Core.scala 44:19]
  assign ifu_io_jump_pc = idu_io_jump_pc; // @[Core.scala 45:19]
  assign ifu_io_en = stall | dmem_not_ok; // @[Core.scala 204:26]
  assign ifu_io_pc = idreg_io_pc_out; // @[Core.scala 46:19]
  assign idu_io_pc = idreg_io_pc_out; // @[Core.scala 54:19]
  assign idu_io_inst = idreg_io_inst_out; // @[Core.scala 55:19]
  assign idu_io_rs1_data = rfu_io_rs1_data; // @[Core.scala 56:19]
  assign idu_io_rs2_data = rfu_io_rs2_data; // @[Core.scala 57:19]
  assign idu_io_mtvec = csru_io_mtvec; // @[Core.scala 58:19]
  assign idu_io_mepc = csru_io_mepc; // @[Core.scala 59:19]
  assign ieu_io_decode_info_alu_code = exereg_io_decode_info_out_alu_code; // @[Core.scala 72:22]
  assign ieu_io_decode_info_bu_code = exereg_io_decode_info_out_bu_code; // @[Core.scala 72:22]
  assign ieu_io_decode_info_mdu_code = exereg_io_decode_info_out_mdu_code; // @[Core.scala 72:22]
  assign ieu_io_decode_info_csru_code = exereg_io_decode_info_out_csru_code; // @[Core.scala 72:22]
  assign ieu_io_op1 = exereg_io_op1_out; // @[Core.scala 73:14]
  assign ieu_io_op2 = exereg_io_op2_out; // @[Core.scala 74:14]
  assign ieu_io_pc = exereg_io_pc_out; // @[Core.scala 75:14]
  assign ieu_io_rs1_addr = exereg_io_rs1_addr_out; // @[Core.scala 77:19]
  assign ieu_io_csr_rdata = csru_io_rdata; // @[Core.scala 79:20]
  assign rfu_clock = clock;
  assign rfu_reset = reset;
  assign rfu_io_rs1_addr = idu_io_rs1_addr; // @[Core.scala 146:19]
  assign rfu_io_rs2_addr = idu_io_rs2_addr; // @[Core.scala 147:19]
  assign rfu_io_rd_addr = wbreg_io_rd_addr_out; // @[Core.scala 149:19]
  assign rfu_io_rd_data = wbu_io_out; // @[Core.scala 151:19]
  assign rfu_io_rd_en = wbreg_io_rd_en_out & commit_valid; // @[Core.scala 205:39]
  assign csru_clock = clock;
  assign csru_reset = reset;
  assign csru_io_raddr = ieu_io_csr_raddr; // @[Core.scala 154:21]
  assign csru_io_wen = wbreg_io_csr_wen_out & commit_valid; // @[Core.scala 206:41]
  assign csru_io_waddr = wbreg_io_csr_waddr_out; // @[Core.scala 155:21]
  assign csru_io_wdata = wbreg_io_csr_wdata_out; // @[Core.scala 156:21]
  assign csru_io_csru_code_valid = wbreg_io_pr_valid_out & ~dmem_not_ok; // @[Core.scala 196:44]
  assign csru_io_csru_code = wbreg_io_csru_code_out; // @[Core.scala 157:21]
  assign csru_io_pc = wbreg_io_pc_out; // @[Core.scala 158:21]
  assign preamu_io_lu_code = memreg_io_decode_info_out_lu_code; // @[Core.scala 100:21]
  assign preamu_io_su_code = memreg_io_decode_info_out_su_code; // @[Core.scala 101:21]
  assign preamu_io_op1 = memreg_io_op1_out; // @[Core.scala 102:21]
  assign preamu_io_op2 = memreg_io_op2_out; // @[Core.scala 103:21]
  assign preamu_io_imm = memreg_io_imm_out; // @[Core.scala 104:21]
  assign amu_io_lu_code = wbreg_io_lu_code_out; // @[Core.scala 134:19]
  assign amu_io_lu_shift = wbreg_io_lu_shift_out; // @[Core.scala 135:19]
  assign amu_io_rdata = io_dmem_rdata; // @[Core.scala 136:19]
  assign wbu_io_fu_code = wbreg_io_fu_code_out; // @[Core.scala 138:19]
  assign wbu_io_alu_out = wbreg_io_alu_out_out; // @[Core.scala 139:19]
  assign wbu_io_bu_out = wbreg_io_bu_out_out; // @[Core.scala 140:19]
  assign wbu_io_mdu_out = wbreg_io_mdu_out_out; // @[Core.scala 141:19]
  assign wbu_io_lu_out = amu_io_lu_out; // @[Core.scala 143:19]
  assign wbu_io_csru_out = wbreg_io_csru_out_out; // @[Core.scala 142:19]
  assign rfconflict_io_rs_valid = idreg_io_pr_valid_out; // @[Core.scala 162:29]
  assign rfconflict_io_rs1_en = idu_io_rs1_en; // @[Core.scala 163:28]
  assign rfconflict_io_rs2_en = idu_io_rs2_en; // @[Core.scala 164:28]
  assign rfconflict_io_rs1_addr = idu_io_rs1_addr; // @[Core.scala 165:28]
  assign rfconflict_io_rs2_addr = idu_io_rs2_addr; // @[Core.scala 166:28]
  assign rfconflict_io_rd1_valid = exereg_io_pr_valid_out; // @[Core.scala 167:28]
  assign rfconflict_io_rd1_en = exereg_io_rd_en_out; // @[Core.scala 168:28]
  assign rfconflict_io_rd1_addr = exereg_io_rd_addr_out; // @[Core.scala 169:28]
  assign rfconflict_io_rd2_valid = memreg_io_pr_valid_out; // @[Core.scala 170:28]
  assign rfconflict_io_rd2_en = memreg_io_rd_en_out; // @[Core.scala 171:28]
  assign rfconflict_io_rd2_addr = memreg_io_rd_addr_out; // @[Core.scala 172:28]
  assign rfconflict_io_rd3_valid = wbreg_io_pr_valid_out; // @[Core.scala 173:28]
  assign rfconflict_io_rd3_en = wbreg_io_rd_en_out; // @[Core.scala 174:28]
  assign rfconflict_io_rd3_addr = wbreg_io_rd_addr_out; // @[Core.scala 175:28]
  assign idreg_clock = clock;
  assign idreg_reset = reset;
  assign idreg_io_imem_data = io_imem_data; // @[Core.scala 50:23]
  assign idreg_io_pr_valid_in = ifu_io_valid; // @[Core.scala 192:25]
  assign idreg_io_pr_en = _exereg_io_pr_valid_in_T & _commit_valid_T; // @[Core.scala 198:29]
  assign idreg_io_pc_in = ifu_io_next_pc; // @[Core.scala 52:19]
  assign exereg_clock = clock;
  assign exereg_reset = reset;
  assign exereg_io_pr_valid_in = idreg_io_pr_valid_out & ~stall; // @[Core.scala 193:50]
  assign exereg_io_pr_en = ~dmem_not_ok; // @[Core.scala 199:22]
  assign exereg_io_pc_in = idreg_io_pc_out; // @[Core.scala 61:25]
  assign exereg_io_inst_in = idreg_io_inst_out; // @[Core.scala 62:25]
  assign exereg_io_rd_en_in = idu_io_rd_en; // @[Core.scala 63:25]
  assign exereg_io_rd_addr_in = idu_io_rd_addr; // @[Core.scala 64:25]
  assign exereg_io_imm_in = idu_io_imm; // @[Core.scala 65:25]
  assign exereg_io_op1_in = idu_io_op1; // @[Core.scala 66:25]
  assign exereg_io_op2_in = idu_io_op2; // @[Core.scala 67:25]
  assign exereg_io_rs1_addr_in = idu_io_rs1_addr; // @[Core.scala 68:25]
  assign exereg_io_decode_info_in_fu_code = idu_io_decode_info_fu_code; // @[Core.scala 69:28]
  assign exereg_io_decode_info_in_alu_code = idu_io_decode_info_alu_code; // @[Core.scala 69:28]
  assign exereg_io_decode_info_in_bu_code = idu_io_decode_info_bu_code; // @[Core.scala 69:28]
  assign exereg_io_decode_info_in_lu_code = idu_io_decode_info_lu_code; // @[Core.scala 69:28]
  assign exereg_io_decode_info_in_su_code = idu_io_decode_info_su_code; // @[Core.scala 69:28]
  assign exereg_io_decode_info_in_mdu_code = idu_io_decode_info_mdu_code; // @[Core.scala 69:28]
  assign exereg_io_decode_info_in_csru_code = idu_io_decode_info_csru_code; // @[Core.scala 69:28]
  assign exereg_io_putch_in = idu_io_putch; // @[Core.scala 70:25]
  assign memreg_clock = clock;
  assign memreg_reset = reset;
  assign memreg_io_pr_valid_in = exereg_io_pr_valid_out; // @[Core.scala 194:25]
  assign memreg_io_pr_en = ~dmem_not_ok; // @[Core.scala 200:22]
  assign memreg_io_pc_in = exereg_io_pc_out; // @[Core.scala 81:25]
  assign memreg_io_inst_in = exereg_io_inst_out; // @[Core.scala 82:25]
  assign memreg_io_rd_en_in = exereg_io_rd_en_out; // @[Core.scala 83:25]
  assign memreg_io_rd_addr_in = exereg_io_rd_addr_out; // @[Core.scala 84:25]
  assign memreg_io_alu_out_in = ieu_io_alu_out; // @[Core.scala 90:25]
  assign memreg_io_bu_out_in = ieu_io_bu_out; // @[Core.scala 91:25]
  assign memreg_io_mdu_out_in = ieu_io_mdu_out; // @[Core.scala 92:25]
  assign memreg_io_csru_out_in = ieu_io_csru_out; // @[Core.scala 93:25]
  assign memreg_io_imm_in = exereg_io_imm_out; // @[Core.scala 85:25]
  assign memreg_io_op1_in = exereg_io_op1_out; // @[Core.scala 86:25]
  assign memreg_io_op2_in = exereg_io_op2_out; // @[Core.scala 87:25]
  assign memreg_io_decode_info_in_fu_code = exereg_io_decode_info_out_fu_code; // @[Core.scala 88:28]
  assign memreg_io_decode_info_in_lu_code = exereg_io_decode_info_out_lu_code; // @[Core.scala 88:28]
  assign memreg_io_decode_info_in_su_code = exereg_io_decode_info_out_su_code; // @[Core.scala 88:28]
  assign memreg_io_decode_info_in_csru_code = exereg_io_decode_info_out_csru_code; // @[Core.scala 88:28]
  assign memreg_io_putch_in = exereg_io_putch_out; // @[Core.scala 95:27]
  assign memreg_io_csr_wen_in = ieu_io_csr_wen; // @[Core.scala 96:27]
  assign memreg_io_csr_waddr_in = ieu_io_csr_waddr; // @[Core.scala 97:27]
  assign memreg_io_csr_wdata_in = ieu_io_csr_wdata; // @[Core.scala 98:27]
  assign wbreg_clock = clock;
  assign wbreg_reset = reset;
  assign wbreg_io_pr_valid_in = memreg_io_pr_valid_out; // @[Core.scala 195:25]
  assign wbreg_io_pr_en = ~dmem_not_ok; // @[Core.scala 201:22]
  assign wbreg_io_pc_in = memreg_io_pc_out; // @[Core.scala 115:25]
  assign wbreg_io_inst_in = memreg_io_inst_out; // @[Core.scala 116:25]
  assign wbreg_io_rd_en_in = memreg_io_rd_en_out; // @[Core.scala 117:25]
  assign wbreg_io_rd_addr_in = memreg_io_rd_addr_out; // @[Core.scala 118:25]
  assign wbreg_io_alu_out_in = memreg_io_alu_out_out; // @[Core.scala 119:25]
  assign wbreg_io_bu_out_in = memreg_io_bu_out_out; // @[Core.scala 120:25]
  assign wbreg_io_mdu_out_in = memreg_io_mdu_out_out; // @[Core.scala 121:25]
  assign wbreg_io_csru_out_in = memreg_io_csru_out_out; // @[Core.scala 122:25]
  assign wbreg_io_fu_code_in = memreg_io_decode_info_out_fu_code; // @[Core.scala 123:25]
  assign wbreg_io_lu_code_in = memreg_io_decode_info_out_lu_code; // @[Core.scala 124:25]
  assign wbreg_io_csru_code_in = memreg_io_decode_info_out_csru_code; // @[Core.scala 125:25]
  assign wbreg_io_lu_shift_in = preamu_io_lu_shift; // @[Core.scala 127:24]
  assign wbreg_io_putch_in = memreg_io_putch_out; // @[Core.scala 129:25]
  assign wbreg_io_csr_wen_in = memreg_io_csr_wen_out; // @[Core.scala 130:25]
  assign wbreg_io_csr_waddr_in = memreg_io_csr_waddr_out; // @[Core.scala 131:25]
  assign wbreg_io_csr_wdata_in = memreg_io_csr_wdata_out; // @[Core.scala 132:25]
  assign dt_ic_clock = clock; // @[Core.scala 225:21]
  assign dt_ic_coreid = 8'h0; // @[Core.scala 226:21]
  assign dt_ic_index = 8'h0; // @[Core.scala 227:21]
  assign dt_ic_valid = dt_ic_io_valid_REG; // @[Core.scala 228:21]
  assign dt_ic_pc = dt_ic_io_pc_REG; // @[Core.scala 229:21]
  assign dt_ic_instr = dt_ic_io_instr_REG; // @[Core.scala 230:21]
  assign dt_ic_special = 8'h0; // @[Core.scala 231:21]
  assign dt_ic_skip = dt_ic_io_skip_REG; // @[Core.scala 232:21]
  assign dt_ic_isRVC = 1'h0; // @[Core.scala 233:21]
  assign dt_ic_scFailed = 1'h0; // @[Core.scala 234:21]
  assign dt_ic_wen = dt_ic_io_wen_REG; // @[Core.scala 235:21]
  assign dt_ic_wdata = dt_ic_io_wdata_REG; // @[Core.scala 236:21]
  assign dt_ic_wdest = {{3'd0}, dt_ic_io_wdest_REG}; // @[Core.scala 237:21]
  assign dt_ae_clock = clock; // @[Core.scala 240:25]
  assign dt_ae_coreid = 8'h0; // @[Core.scala 241:25]
  assign dt_ae_intrNO = 32'h0; // @[Core.scala 242:25]
  assign dt_ae_cause = 32'h0; // @[Core.scala 243:25]
  assign dt_ae_exceptionPC = 64'h0; // @[Core.scala 244:25]
  assign dt_ae_exceptionInst = 32'h0;
  assign dt_te_clock = clock; // @[Core.scala 256:21]
  assign dt_te_coreid = 8'h0; // @[Core.scala 257:21]
  assign dt_te_valid = wbreg_io_inst_out == 32'h6b & commit_valid; // @[Core.scala 258:62]
  assign dt_te_code = rf_a0_0[2:0]; // @[Core.scala 259:29]
  assign dt_te_pc = wbreg_io_pc_out; // @[Core.scala 260:21]
  assign dt_te_cycleCnt = cycle_cnt; // @[Core.scala 261:21]
  assign dt_te_instrCnt = instr_cnt; // @[Core.scala 262:21]
  always @(posedge clock) begin
    dt_ic_io_valid_REG <= wbreg_io_pr_valid_out & ~dmem_not_ok; // @[Core.scala 196:44]
    dt_ic_io_pc_REG <= wbreg_io_pc_out; // @[Core.scala 229:31]
    dt_ic_io_instr_REG <= wbreg_io_inst_out; // @[Core.scala 230:31]
    dt_ic_io_skip_REG <= wbreg_io_inst_out == 32'h7b | read_mcycle | read_mtime | write_mtimecmp | wbreg_io_inst_out == 32'h7b703
      ; // @[Core.scala 232:107]
    dt_ic_io_wen_REG <= wbreg_io_rd_en_out; // @[Core.scala 235:31]
    dt_ic_io_wdata_REG <= wbu_io_out; // @[Core.scala 236:31]
    dt_ic_io_wdest_REG <= wbreg_io_rd_addr_out; // @[Core.scala 237:31]
    if (reset) begin // @[Core.scala 246:26]
      cycle_cnt <= 64'h0; // @[Core.scala 246:26]
    end else begin
      cycle_cnt <= _cycle_cnt_T_1; // @[Core.scala 249:13]
    end
    if (reset) begin // @[Core.scala 247:26]
      instr_cnt <= 64'h0; // @[Core.scala 247:26]
    end else if (commit_valid) begin // @[Core.scala 250:19]
      instr_cnt <= _instr_cnt_T_1;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (wbreg_io_putch_out & commit_valid & ~reset) begin
          $fwrite(32'h80000002,"%c",rf_a0_0); // @[Core.scala 213:51]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  dt_ic_io_valid_REG = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  dt_ic_io_pc_REG = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  dt_ic_io_instr_REG = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  dt_ic_io_skip_REG = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  dt_ic_io_wen_REG = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  dt_ic_io_wdata_REG = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  dt_ic_io_wdest_REG = _RAND_6[4:0];
  _RAND_7 = {2{`RANDOM}};
  cycle_cnt = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  instr_cnt = _RAND_8[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ICache(
  input          clock,
  input          reset,
  input  [63:0]  io_imem_addr,
  output [31:0]  io_imem_data,
  output         io_imem_data_ok,
  output         io_axi_req,
  output [63:0]  io_axi_addr,
  input          io_axi_valid,
  input  [511:0] io_axi_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [63:0] _RAND_65;
  reg [63:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [63:0] _RAND_68;
  reg [63:0] _RAND_69;
  reg [63:0] _RAND_70;
  reg [63:0] _RAND_71;
  reg [63:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [63:0] _RAND_75;
  reg [63:0] _RAND_76;
  reg [63:0] _RAND_77;
  reg [63:0] _RAND_78;
  reg [63:0] _RAND_79;
  reg [63:0] _RAND_80;
  reg [63:0] _RAND_81;
  reg [63:0] _RAND_82;
  reg [63:0] _RAND_83;
  reg [63:0] _RAND_84;
  reg [63:0] _RAND_85;
  reg [63:0] _RAND_86;
  reg [63:0] _RAND_87;
  reg [63:0] _RAND_88;
  reg [63:0] _RAND_89;
  reg [63:0] _RAND_90;
  reg [63:0] _RAND_91;
  reg [63:0] _RAND_92;
  reg [63:0] _RAND_93;
  reg [63:0] _RAND_94;
  reg [63:0] _RAND_95;
  reg [511:0] _RAND_96;
  reg [511:0] _RAND_97;
  reg [511:0] _RAND_98;
  reg [511:0] _RAND_99;
  reg [511:0] _RAND_100;
  reg [511:0] _RAND_101;
  reg [511:0] _RAND_102;
  reg [511:0] _RAND_103;
  reg [511:0] _RAND_104;
  reg [511:0] _RAND_105;
  reg [511:0] _RAND_106;
  reg [511:0] _RAND_107;
  reg [511:0] _RAND_108;
  reg [511:0] _RAND_109;
  reg [511:0] _RAND_110;
  reg [511:0] _RAND_111;
  reg [511:0] _RAND_112;
  reg [511:0] _RAND_113;
  reg [511:0] _RAND_114;
  reg [511:0] _RAND_115;
  reg [511:0] _RAND_116;
  reg [511:0] _RAND_117;
  reg [511:0] _RAND_118;
  reg [511:0] _RAND_119;
  reg [511:0] _RAND_120;
  reg [511:0] _RAND_121;
  reg [511:0] _RAND_122;
  reg [511:0] _RAND_123;
  reg [511:0] _RAND_124;
  reg [511:0] _RAND_125;
  reg [511:0] _RAND_126;
  reg [511:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [63:0] _RAND_192;
  reg [63:0] _RAND_193;
  reg [63:0] _RAND_194;
  reg [63:0] _RAND_195;
  reg [63:0] _RAND_196;
  reg [63:0] _RAND_197;
  reg [63:0] _RAND_198;
  reg [63:0] _RAND_199;
  reg [63:0] _RAND_200;
  reg [63:0] _RAND_201;
  reg [63:0] _RAND_202;
  reg [63:0] _RAND_203;
  reg [63:0] _RAND_204;
  reg [63:0] _RAND_205;
  reg [63:0] _RAND_206;
  reg [63:0] _RAND_207;
  reg [63:0] _RAND_208;
  reg [63:0] _RAND_209;
  reg [63:0] _RAND_210;
  reg [63:0] _RAND_211;
  reg [63:0] _RAND_212;
  reg [63:0] _RAND_213;
  reg [63:0] _RAND_214;
  reg [63:0] _RAND_215;
  reg [63:0] _RAND_216;
  reg [63:0] _RAND_217;
  reg [63:0] _RAND_218;
  reg [63:0] _RAND_219;
  reg [63:0] _RAND_220;
  reg [63:0] _RAND_221;
  reg [63:0] _RAND_222;
  reg [63:0] _RAND_223;
  reg [511:0] _RAND_224;
  reg [511:0] _RAND_225;
  reg [511:0] _RAND_226;
  reg [511:0] _RAND_227;
  reg [511:0] _RAND_228;
  reg [511:0] _RAND_229;
  reg [511:0] _RAND_230;
  reg [511:0] _RAND_231;
  reg [511:0] _RAND_232;
  reg [511:0] _RAND_233;
  reg [511:0] _RAND_234;
  reg [511:0] _RAND_235;
  reg [511:0] _RAND_236;
  reg [511:0] _RAND_237;
  reg [511:0] _RAND_238;
  reg [511:0] _RAND_239;
  reg [511:0] _RAND_240;
  reg [511:0] _RAND_241;
  reg [511:0] _RAND_242;
  reg [511:0] _RAND_243;
  reg [511:0] _RAND_244;
  reg [511:0] _RAND_245;
  reg [511:0] _RAND_246;
  reg [511:0] _RAND_247;
  reg [511:0] _RAND_248;
  reg [511:0] _RAND_249;
  reg [511:0] _RAND_250;
  reg [511:0] _RAND_251;
  reg [511:0] _RAND_252;
  reg [511:0] _RAND_253;
  reg [511:0] _RAND_254;
  reg [511:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
`endif // RANDOMIZE_REG_INIT
  wire [52:0] tag_addr = io_imem_addr[63:11]; // @[ICache.scala 43:35]
  wire [4:0] index_addr = io_imem_addr[10:6]; // @[ICache.scala 44:35]
  wire [5:0] offset_addr = io_imem_addr[5:0]; // @[ICache.scala 45:35]
  reg  v1_0; // @[ICache.scala 47:26]
  reg  v1_1; // @[ICache.scala 47:26]
  reg  v1_2; // @[ICache.scala 47:26]
  reg  v1_3; // @[ICache.scala 47:26]
  reg  v1_4; // @[ICache.scala 47:26]
  reg  v1_5; // @[ICache.scala 47:26]
  reg  v1_6; // @[ICache.scala 47:26]
  reg  v1_7; // @[ICache.scala 47:26]
  reg  v1_8; // @[ICache.scala 47:26]
  reg  v1_9; // @[ICache.scala 47:26]
  reg  v1_10; // @[ICache.scala 47:26]
  reg  v1_11; // @[ICache.scala 47:26]
  reg  v1_12; // @[ICache.scala 47:26]
  reg  v1_13; // @[ICache.scala 47:26]
  reg  v1_14; // @[ICache.scala 47:26]
  reg  v1_15; // @[ICache.scala 47:26]
  reg  v1_16; // @[ICache.scala 47:26]
  reg  v1_17; // @[ICache.scala 47:26]
  reg  v1_18; // @[ICache.scala 47:26]
  reg  v1_19; // @[ICache.scala 47:26]
  reg  v1_20; // @[ICache.scala 47:26]
  reg  v1_21; // @[ICache.scala 47:26]
  reg  v1_22; // @[ICache.scala 47:26]
  reg  v1_23; // @[ICache.scala 47:26]
  reg  v1_24; // @[ICache.scala 47:26]
  reg  v1_25; // @[ICache.scala 47:26]
  reg  v1_26; // @[ICache.scala 47:26]
  reg  v1_27; // @[ICache.scala 47:26]
  reg  v1_28; // @[ICache.scala 47:26]
  reg  v1_29; // @[ICache.scala 47:26]
  reg  v1_30; // @[ICache.scala 47:26]
  reg  v1_31; // @[ICache.scala 47:26]
  reg  age1_0; // @[ICache.scala 48:26]
  reg  age1_1; // @[ICache.scala 48:26]
  reg  age1_2; // @[ICache.scala 48:26]
  reg  age1_3; // @[ICache.scala 48:26]
  reg  age1_4; // @[ICache.scala 48:26]
  reg  age1_5; // @[ICache.scala 48:26]
  reg  age1_6; // @[ICache.scala 48:26]
  reg  age1_7; // @[ICache.scala 48:26]
  reg  age1_8; // @[ICache.scala 48:26]
  reg  age1_9; // @[ICache.scala 48:26]
  reg  age1_10; // @[ICache.scala 48:26]
  reg  age1_11; // @[ICache.scala 48:26]
  reg  age1_12; // @[ICache.scala 48:26]
  reg  age1_13; // @[ICache.scala 48:26]
  reg  age1_14; // @[ICache.scala 48:26]
  reg  age1_15; // @[ICache.scala 48:26]
  reg  age1_16; // @[ICache.scala 48:26]
  reg  age1_17; // @[ICache.scala 48:26]
  reg  age1_18; // @[ICache.scala 48:26]
  reg  age1_19; // @[ICache.scala 48:26]
  reg  age1_20; // @[ICache.scala 48:26]
  reg  age1_21; // @[ICache.scala 48:26]
  reg  age1_22; // @[ICache.scala 48:26]
  reg  age1_23; // @[ICache.scala 48:26]
  reg  age1_24; // @[ICache.scala 48:26]
  reg  age1_25; // @[ICache.scala 48:26]
  reg  age1_26; // @[ICache.scala 48:26]
  reg  age1_27; // @[ICache.scala 48:26]
  reg  age1_28; // @[ICache.scala 48:26]
  reg  age1_29; // @[ICache.scala 48:26]
  reg  age1_30; // @[ICache.scala 48:26]
  reg  age1_31; // @[ICache.scala 48:26]
  reg [52:0] tag1_0; // @[ICache.scala 49:26]
  reg [52:0] tag1_1; // @[ICache.scala 49:26]
  reg [52:0] tag1_2; // @[ICache.scala 49:26]
  reg [52:0] tag1_3; // @[ICache.scala 49:26]
  reg [52:0] tag1_4; // @[ICache.scala 49:26]
  reg [52:0] tag1_5; // @[ICache.scala 49:26]
  reg [52:0] tag1_6; // @[ICache.scala 49:26]
  reg [52:0] tag1_7; // @[ICache.scala 49:26]
  reg [52:0] tag1_8; // @[ICache.scala 49:26]
  reg [52:0] tag1_9; // @[ICache.scala 49:26]
  reg [52:0] tag1_10; // @[ICache.scala 49:26]
  reg [52:0] tag1_11; // @[ICache.scala 49:26]
  reg [52:0] tag1_12; // @[ICache.scala 49:26]
  reg [52:0] tag1_13; // @[ICache.scala 49:26]
  reg [52:0] tag1_14; // @[ICache.scala 49:26]
  reg [52:0] tag1_15; // @[ICache.scala 49:26]
  reg [52:0] tag1_16; // @[ICache.scala 49:26]
  reg [52:0] tag1_17; // @[ICache.scala 49:26]
  reg [52:0] tag1_18; // @[ICache.scala 49:26]
  reg [52:0] tag1_19; // @[ICache.scala 49:26]
  reg [52:0] tag1_20; // @[ICache.scala 49:26]
  reg [52:0] tag1_21; // @[ICache.scala 49:26]
  reg [52:0] tag1_22; // @[ICache.scala 49:26]
  reg [52:0] tag1_23; // @[ICache.scala 49:26]
  reg [52:0] tag1_24; // @[ICache.scala 49:26]
  reg [52:0] tag1_25; // @[ICache.scala 49:26]
  reg [52:0] tag1_26; // @[ICache.scala 49:26]
  reg [52:0] tag1_27; // @[ICache.scala 49:26]
  reg [52:0] tag1_28; // @[ICache.scala 49:26]
  reg [52:0] tag1_29; // @[ICache.scala 49:26]
  reg [52:0] tag1_30; // @[ICache.scala 49:26]
  reg [52:0] tag1_31; // @[ICache.scala 49:26]
  reg [511:0] block1_0; // @[ICache.scala 50:26]
  reg [511:0] block1_1; // @[ICache.scala 50:26]
  reg [511:0] block1_2; // @[ICache.scala 50:26]
  reg [511:0] block1_3; // @[ICache.scala 50:26]
  reg [511:0] block1_4; // @[ICache.scala 50:26]
  reg [511:0] block1_5; // @[ICache.scala 50:26]
  reg [511:0] block1_6; // @[ICache.scala 50:26]
  reg [511:0] block1_7; // @[ICache.scala 50:26]
  reg [511:0] block1_8; // @[ICache.scala 50:26]
  reg [511:0] block1_9; // @[ICache.scala 50:26]
  reg [511:0] block1_10; // @[ICache.scala 50:26]
  reg [511:0] block1_11; // @[ICache.scala 50:26]
  reg [511:0] block1_12; // @[ICache.scala 50:26]
  reg [511:0] block1_13; // @[ICache.scala 50:26]
  reg [511:0] block1_14; // @[ICache.scala 50:26]
  reg [511:0] block1_15; // @[ICache.scala 50:26]
  reg [511:0] block1_16; // @[ICache.scala 50:26]
  reg [511:0] block1_17; // @[ICache.scala 50:26]
  reg [511:0] block1_18; // @[ICache.scala 50:26]
  reg [511:0] block1_19; // @[ICache.scala 50:26]
  reg [511:0] block1_20; // @[ICache.scala 50:26]
  reg [511:0] block1_21; // @[ICache.scala 50:26]
  reg [511:0] block1_22; // @[ICache.scala 50:26]
  reg [511:0] block1_23; // @[ICache.scala 50:26]
  reg [511:0] block1_24; // @[ICache.scala 50:26]
  reg [511:0] block1_25; // @[ICache.scala 50:26]
  reg [511:0] block1_26; // @[ICache.scala 50:26]
  reg [511:0] block1_27; // @[ICache.scala 50:26]
  reg [511:0] block1_28; // @[ICache.scala 50:26]
  reg [511:0] block1_29; // @[ICache.scala 50:26]
  reg [511:0] block1_30; // @[ICache.scala 50:26]
  reg [511:0] block1_31; // @[ICache.scala 50:26]
  reg  v2_0; // @[ICache.scala 51:26]
  reg  v2_1; // @[ICache.scala 51:26]
  reg  v2_2; // @[ICache.scala 51:26]
  reg  v2_3; // @[ICache.scala 51:26]
  reg  v2_4; // @[ICache.scala 51:26]
  reg  v2_5; // @[ICache.scala 51:26]
  reg  v2_6; // @[ICache.scala 51:26]
  reg  v2_7; // @[ICache.scala 51:26]
  reg  v2_8; // @[ICache.scala 51:26]
  reg  v2_9; // @[ICache.scala 51:26]
  reg  v2_10; // @[ICache.scala 51:26]
  reg  v2_11; // @[ICache.scala 51:26]
  reg  v2_12; // @[ICache.scala 51:26]
  reg  v2_13; // @[ICache.scala 51:26]
  reg  v2_14; // @[ICache.scala 51:26]
  reg  v2_15; // @[ICache.scala 51:26]
  reg  v2_16; // @[ICache.scala 51:26]
  reg  v2_17; // @[ICache.scala 51:26]
  reg  v2_18; // @[ICache.scala 51:26]
  reg  v2_19; // @[ICache.scala 51:26]
  reg  v2_20; // @[ICache.scala 51:26]
  reg  v2_21; // @[ICache.scala 51:26]
  reg  v2_22; // @[ICache.scala 51:26]
  reg  v2_23; // @[ICache.scala 51:26]
  reg  v2_24; // @[ICache.scala 51:26]
  reg  v2_25; // @[ICache.scala 51:26]
  reg  v2_26; // @[ICache.scala 51:26]
  reg  v2_27; // @[ICache.scala 51:26]
  reg  v2_28; // @[ICache.scala 51:26]
  reg  v2_29; // @[ICache.scala 51:26]
  reg  v2_30; // @[ICache.scala 51:26]
  reg  v2_31; // @[ICache.scala 51:26]
  reg  age2_0; // @[ICache.scala 52:26]
  reg  age2_1; // @[ICache.scala 52:26]
  reg  age2_2; // @[ICache.scala 52:26]
  reg  age2_3; // @[ICache.scala 52:26]
  reg  age2_4; // @[ICache.scala 52:26]
  reg  age2_5; // @[ICache.scala 52:26]
  reg  age2_6; // @[ICache.scala 52:26]
  reg  age2_7; // @[ICache.scala 52:26]
  reg  age2_8; // @[ICache.scala 52:26]
  reg  age2_9; // @[ICache.scala 52:26]
  reg  age2_10; // @[ICache.scala 52:26]
  reg  age2_11; // @[ICache.scala 52:26]
  reg  age2_12; // @[ICache.scala 52:26]
  reg  age2_13; // @[ICache.scala 52:26]
  reg  age2_14; // @[ICache.scala 52:26]
  reg  age2_15; // @[ICache.scala 52:26]
  reg  age2_16; // @[ICache.scala 52:26]
  reg  age2_17; // @[ICache.scala 52:26]
  reg  age2_18; // @[ICache.scala 52:26]
  reg  age2_19; // @[ICache.scala 52:26]
  reg  age2_20; // @[ICache.scala 52:26]
  reg  age2_21; // @[ICache.scala 52:26]
  reg  age2_22; // @[ICache.scala 52:26]
  reg  age2_23; // @[ICache.scala 52:26]
  reg  age2_24; // @[ICache.scala 52:26]
  reg  age2_25; // @[ICache.scala 52:26]
  reg  age2_26; // @[ICache.scala 52:26]
  reg  age2_27; // @[ICache.scala 52:26]
  reg  age2_28; // @[ICache.scala 52:26]
  reg  age2_29; // @[ICache.scala 52:26]
  reg  age2_30; // @[ICache.scala 52:26]
  reg  age2_31; // @[ICache.scala 52:26]
  reg [52:0] tag2_0; // @[ICache.scala 53:26]
  reg [52:0] tag2_1; // @[ICache.scala 53:26]
  reg [52:0] tag2_2; // @[ICache.scala 53:26]
  reg [52:0] tag2_3; // @[ICache.scala 53:26]
  reg [52:0] tag2_4; // @[ICache.scala 53:26]
  reg [52:0] tag2_5; // @[ICache.scala 53:26]
  reg [52:0] tag2_6; // @[ICache.scala 53:26]
  reg [52:0] tag2_7; // @[ICache.scala 53:26]
  reg [52:0] tag2_8; // @[ICache.scala 53:26]
  reg [52:0] tag2_9; // @[ICache.scala 53:26]
  reg [52:0] tag2_10; // @[ICache.scala 53:26]
  reg [52:0] tag2_11; // @[ICache.scala 53:26]
  reg [52:0] tag2_12; // @[ICache.scala 53:26]
  reg [52:0] tag2_13; // @[ICache.scala 53:26]
  reg [52:0] tag2_14; // @[ICache.scala 53:26]
  reg [52:0] tag2_15; // @[ICache.scala 53:26]
  reg [52:0] tag2_16; // @[ICache.scala 53:26]
  reg [52:0] tag2_17; // @[ICache.scala 53:26]
  reg [52:0] tag2_18; // @[ICache.scala 53:26]
  reg [52:0] tag2_19; // @[ICache.scala 53:26]
  reg [52:0] tag2_20; // @[ICache.scala 53:26]
  reg [52:0] tag2_21; // @[ICache.scala 53:26]
  reg [52:0] tag2_22; // @[ICache.scala 53:26]
  reg [52:0] tag2_23; // @[ICache.scala 53:26]
  reg [52:0] tag2_24; // @[ICache.scala 53:26]
  reg [52:0] tag2_25; // @[ICache.scala 53:26]
  reg [52:0] tag2_26; // @[ICache.scala 53:26]
  reg [52:0] tag2_27; // @[ICache.scala 53:26]
  reg [52:0] tag2_28; // @[ICache.scala 53:26]
  reg [52:0] tag2_29; // @[ICache.scala 53:26]
  reg [52:0] tag2_30; // @[ICache.scala 53:26]
  reg [52:0] tag2_31; // @[ICache.scala 53:26]
  reg [511:0] block2_0; // @[ICache.scala 54:26]
  reg [511:0] block2_1; // @[ICache.scala 54:26]
  reg [511:0] block2_2; // @[ICache.scala 54:26]
  reg [511:0] block2_3; // @[ICache.scala 54:26]
  reg [511:0] block2_4; // @[ICache.scala 54:26]
  reg [511:0] block2_5; // @[ICache.scala 54:26]
  reg [511:0] block2_6; // @[ICache.scala 54:26]
  reg [511:0] block2_7; // @[ICache.scala 54:26]
  reg [511:0] block2_8; // @[ICache.scala 54:26]
  reg [511:0] block2_9; // @[ICache.scala 54:26]
  reg [511:0] block2_10; // @[ICache.scala 54:26]
  reg [511:0] block2_11; // @[ICache.scala 54:26]
  reg [511:0] block2_12; // @[ICache.scala 54:26]
  reg [511:0] block2_13; // @[ICache.scala 54:26]
  reg [511:0] block2_14; // @[ICache.scala 54:26]
  reg [511:0] block2_15; // @[ICache.scala 54:26]
  reg [511:0] block2_16; // @[ICache.scala 54:26]
  reg [511:0] block2_17; // @[ICache.scala 54:26]
  reg [511:0] block2_18; // @[ICache.scala 54:26]
  reg [511:0] block2_19; // @[ICache.scala 54:26]
  reg [511:0] block2_20; // @[ICache.scala 54:26]
  reg [511:0] block2_21; // @[ICache.scala 54:26]
  reg [511:0] block2_22; // @[ICache.scala 54:26]
  reg [511:0] block2_23; // @[ICache.scala 54:26]
  reg [511:0] block2_24; // @[ICache.scala 54:26]
  reg [511:0] block2_25; // @[ICache.scala 54:26]
  reg [511:0] block2_26; // @[ICache.scala 54:26]
  reg [511:0] block2_27; // @[ICache.scala 54:26]
  reg [511:0] block2_28; // @[ICache.scala 54:26]
  reg [511:0] block2_29; // @[ICache.scala 54:26]
  reg [511:0] block2_30; // @[ICache.scala 54:26]
  reg [511:0] block2_31; // @[ICache.scala 54:26]
  wire [52:0] _GEN_1 = 5'h1 == index_addr ? tag1_1 : tag1_0; // @[ICache.scala 56:28 ICache.scala 56:28]
  wire [52:0] _GEN_2 = 5'h2 == index_addr ? tag1_2 : _GEN_1; // @[ICache.scala 56:28 ICache.scala 56:28]
  wire [52:0] _GEN_3 = 5'h3 == index_addr ? tag1_3 : _GEN_2; // @[ICache.scala 56:28 ICache.scala 56:28]
  wire [52:0] _GEN_4 = 5'h4 == index_addr ? tag1_4 : _GEN_3; // @[ICache.scala 56:28 ICache.scala 56:28]
  wire [52:0] _GEN_5 = 5'h5 == index_addr ? tag1_5 : _GEN_4; // @[ICache.scala 56:28 ICache.scala 56:28]
  wire [52:0] _GEN_6 = 5'h6 == index_addr ? tag1_6 : _GEN_5; // @[ICache.scala 56:28 ICache.scala 56:28]
  wire [52:0] _GEN_7 = 5'h7 == index_addr ? tag1_7 : _GEN_6; // @[ICache.scala 56:28 ICache.scala 56:28]
  wire [52:0] _GEN_8 = 5'h8 == index_addr ? tag1_8 : _GEN_7; // @[ICache.scala 56:28 ICache.scala 56:28]
  wire [52:0] _GEN_9 = 5'h9 == index_addr ? tag1_9 : _GEN_8; // @[ICache.scala 56:28 ICache.scala 56:28]
  wire [52:0] _GEN_10 = 5'ha == index_addr ? tag1_10 : _GEN_9; // @[ICache.scala 56:28 ICache.scala 56:28]
  wire [52:0] _GEN_11 = 5'hb == index_addr ? tag1_11 : _GEN_10; // @[ICache.scala 56:28 ICache.scala 56:28]
  wire [52:0] _GEN_12 = 5'hc == index_addr ? tag1_12 : _GEN_11; // @[ICache.scala 56:28 ICache.scala 56:28]
  wire [52:0] _GEN_13 = 5'hd == index_addr ? tag1_13 : _GEN_12; // @[ICache.scala 56:28 ICache.scala 56:28]
  wire [52:0] _GEN_14 = 5'he == index_addr ? tag1_14 : _GEN_13; // @[ICache.scala 56:28 ICache.scala 56:28]
  wire [52:0] _GEN_15 = 5'hf == index_addr ? tag1_15 : _GEN_14; // @[ICache.scala 56:28 ICache.scala 56:28]
  wire [52:0] _GEN_16 = 5'h10 == index_addr ? tag1_16 : _GEN_15; // @[ICache.scala 56:28 ICache.scala 56:28]
  wire [52:0] _GEN_17 = 5'h11 == index_addr ? tag1_17 : _GEN_16; // @[ICache.scala 56:28 ICache.scala 56:28]
  wire [52:0] _GEN_18 = 5'h12 == index_addr ? tag1_18 : _GEN_17; // @[ICache.scala 56:28 ICache.scala 56:28]
  wire [52:0] _GEN_19 = 5'h13 == index_addr ? tag1_19 : _GEN_18; // @[ICache.scala 56:28 ICache.scala 56:28]
  wire [52:0] _GEN_20 = 5'h14 == index_addr ? tag1_20 : _GEN_19; // @[ICache.scala 56:28 ICache.scala 56:28]
  wire [52:0] _GEN_21 = 5'h15 == index_addr ? tag1_21 : _GEN_20; // @[ICache.scala 56:28 ICache.scala 56:28]
  wire [52:0] _GEN_22 = 5'h16 == index_addr ? tag1_22 : _GEN_21; // @[ICache.scala 56:28 ICache.scala 56:28]
  wire [52:0] _GEN_23 = 5'h17 == index_addr ? tag1_23 : _GEN_22; // @[ICache.scala 56:28 ICache.scala 56:28]
  wire [52:0] _GEN_24 = 5'h18 == index_addr ? tag1_24 : _GEN_23; // @[ICache.scala 56:28 ICache.scala 56:28]
  wire [52:0] _GEN_25 = 5'h19 == index_addr ? tag1_25 : _GEN_24; // @[ICache.scala 56:28 ICache.scala 56:28]
  wire [52:0] _GEN_26 = 5'h1a == index_addr ? tag1_26 : _GEN_25; // @[ICache.scala 56:28 ICache.scala 56:28]
  wire [52:0] _GEN_27 = 5'h1b == index_addr ? tag1_27 : _GEN_26; // @[ICache.scala 56:28 ICache.scala 56:28]
  wire [52:0] _GEN_28 = 5'h1c == index_addr ? tag1_28 : _GEN_27; // @[ICache.scala 56:28 ICache.scala 56:28]
  wire [52:0] _GEN_29 = 5'h1d == index_addr ? tag1_29 : _GEN_28; // @[ICache.scala 56:28 ICache.scala 56:28]
  wire [52:0] _GEN_30 = 5'h1e == index_addr ? tag1_30 : _GEN_29; // @[ICache.scala 56:28 ICache.scala 56:28]
  wire [52:0] _GEN_31 = 5'h1f == index_addr ? tag1_31 : _GEN_30; // @[ICache.scala 56:28 ICache.scala 56:28]
  wire  _GEN_33 = 5'h1 == index_addr ? v1_1 : v1_0; // @[ICache.scala 56:67 ICache.scala 56:67]
  wire  _GEN_34 = 5'h2 == index_addr ? v1_2 : _GEN_33; // @[ICache.scala 56:67 ICache.scala 56:67]
  wire  _GEN_35 = 5'h3 == index_addr ? v1_3 : _GEN_34; // @[ICache.scala 56:67 ICache.scala 56:67]
  wire  _GEN_36 = 5'h4 == index_addr ? v1_4 : _GEN_35; // @[ICache.scala 56:67 ICache.scala 56:67]
  wire  _GEN_37 = 5'h5 == index_addr ? v1_5 : _GEN_36; // @[ICache.scala 56:67 ICache.scala 56:67]
  wire  _GEN_38 = 5'h6 == index_addr ? v1_6 : _GEN_37; // @[ICache.scala 56:67 ICache.scala 56:67]
  wire  _GEN_39 = 5'h7 == index_addr ? v1_7 : _GEN_38; // @[ICache.scala 56:67 ICache.scala 56:67]
  wire  _GEN_40 = 5'h8 == index_addr ? v1_8 : _GEN_39; // @[ICache.scala 56:67 ICache.scala 56:67]
  wire  _GEN_41 = 5'h9 == index_addr ? v1_9 : _GEN_40; // @[ICache.scala 56:67 ICache.scala 56:67]
  wire  _GEN_42 = 5'ha == index_addr ? v1_10 : _GEN_41; // @[ICache.scala 56:67 ICache.scala 56:67]
  wire  _GEN_43 = 5'hb == index_addr ? v1_11 : _GEN_42; // @[ICache.scala 56:67 ICache.scala 56:67]
  wire  _GEN_44 = 5'hc == index_addr ? v1_12 : _GEN_43; // @[ICache.scala 56:67 ICache.scala 56:67]
  wire  _GEN_45 = 5'hd == index_addr ? v1_13 : _GEN_44; // @[ICache.scala 56:67 ICache.scala 56:67]
  wire  _GEN_46 = 5'he == index_addr ? v1_14 : _GEN_45; // @[ICache.scala 56:67 ICache.scala 56:67]
  wire  _GEN_47 = 5'hf == index_addr ? v1_15 : _GEN_46; // @[ICache.scala 56:67 ICache.scala 56:67]
  wire  _GEN_48 = 5'h10 == index_addr ? v1_16 : _GEN_47; // @[ICache.scala 56:67 ICache.scala 56:67]
  wire  _GEN_49 = 5'h11 == index_addr ? v1_17 : _GEN_48; // @[ICache.scala 56:67 ICache.scala 56:67]
  wire  _GEN_50 = 5'h12 == index_addr ? v1_18 : _GEN_49; // @[ICache.scala 56:67 ICache.scala 56:67]
  wire  _GEN_51 = 5'h13 == index_addr ? v1_19 : _GEN_50; // @[ICache.scala 56:67 ICache.scala 56:67]
  wire  _GEN_52 = 5'h14 == index_addr ? v1_20 : _GEN_51; // @[ICache.scala 56:67 ICache.scala 56:67]
  wire  _GEN_53 = 5'h15 == index_addr ? v1_21 : _GEN_52; // @[ICache.scala 56:67 ICache.scala 56:67]
  wire  _GEN_54 = 5'h16 == index_addr ? v1_22 : _GEN_53; // @[ICache.scala 56:67 ICache.scala 56:67]
  wire  _GEN_55 = 5'h17 == index_addr ? v1_23 : _GEN_54; // @[ICache.scala 56:67 ICache.scala 56:67]
  wire  _GEN_56 = 5'h18 == index_addr ? v1_24 : _GEN_55; // @[ICache.scala 56:67 ICache.scala 56:67]
  wire  _GEN_57 = 5'h19 == index_addr ? v1_25 : _GEN_56; // @[ICache.scala 56:67 ICache.scala 56:67]
  wire  _GEN_58 = 5'h1a == index_addr ? v1_26 : _GEN_57; // @[ICache.scala 56:67 ICache.scala 56:67]
  wire  _GEN_59 = 5'h1b == index_addr ? v1_27 : _GEN_58; // @[ICache.scala 56:67 ICache.scala 56:67]
  wire  _GEN_60 = 5'h1c == index_addr ? v1_28 : _GEN_59; // @[ICache.scala 56:67 ICache.scala 56:67]
  wire  _GEN_61 = 5'h1d == index_addr ? v1_29 : _GEN_60; // @[ICache.scala 56:67 ICache.scala 56:67]
  wire  _GEN_62 = 5'h1e == index_addr ? v1_30 : _GEN_61; // @[ICache.scala 56:67 ICache.scala 56:67]
  wire  _GEN_63 = 5'h1f == index_addr ? v1_31 : _GEN_62; // @[ICache.scala 56:67 ICache.scala 56:67]
  wire  hit1 = tag_addr == _GEN_31 & _GEN_63; // @[ICache.scala 56:49]
  wire [52:0] _GEN_65 = 5'h1 == index_addr ? tag2_1 : tag2_0; // @[ICache.scala 57:28 ICache.scala 57:28]
  wire [52:0] _GEN_66 = 5'h2 == index_addr ? tag2_2 : _GEN_65; // @[ICache.scala 57:28 ICache.scala 57:28]
  wire [52:0] _GEN_67 = 5'h3 == index_addr ? tag2_3 : _GEN_66; // @[ICache.scala 57:28 ICache.scala 57:28]
  wire [52:0] _GEN_68 = 5'h4 == index_addr ? tag2_4 : _GEN_67; // @[ICache.scala 57:28 ICache.scala 57:28]
  wire [52:0] _GEN_69 = 5'h5 == index_addr ? tag2_5 : _GEN_68; // @[ICache.scala 57:28 ICache.scala 57:28]
  wire [52:0] _GEN_70 = 5'h6 == index_addr ? tag2_6 : _GEN_69; // @[ICache.scala 57:28 ICache.scala 57:28]
  wire [52:0] _GEN_71 = 5'h7 == index_addr ? tag2_7 : _GEN_70; // @[ICache.scala 57:28 ICache.scala 57:28]
  wire [52:0] _GEN_72 = 5'h8 == index_addr ? tag2_8 : _GEN_71; // @[ICache.scala 57:28 ICache.scala 57:28]
  wire [52:0] _GEN_73 = 5'h9 == index_addr ? tag2_9 : _GEN_72; // @[ICache.scala 57:28 ICache.scala 57:28]
  wire [52:0] _GEN_74 = 5'ha == index_addr ? tag2_10 : _GEN_73; // @[ICache.scala 57:28 ICache.scala 57:28]
  wire [52:0] _GEN_75 = 5'hb == index_addr ? tag2_11 : _GEN_74; // @[ICache.scala 57:28 ICache.scala 57:28]
  wire [52:0] _GEN_76 = 5'hc == index_addr ? tag2_12 : _GEN_75; // @[ICache.scala 57:28 ICache.scala 57:28]
  wire [52:0] _GEN_77 = 5'hd == index_addr ? tag2_13 : _GEN_76; // @[ICache.scala 57:28 ICache.scala 57:28]
  wire [52:0] _GEN_78 = 5'he == index_addr ? tag2_14 : _GEN_77; // @[ICache.scala 57:28 ICache.scala 57:28]
  wire [52:0] _GEN_79 = 5'hf == index_addr ? tag2_15 : _GEN_78; // @[ICache.scala 57:28 ICache.scala 57:28]
  wire [52:0] _GEN_80 = 5'h10 == index_addr ? tag2_16 : _GEN_79; // @[ICache.scala 57:28 ICache.scala 57:28]
  wire [52:0] _GEN_81 = 5'h11 == index_addr ? tag2_17 : _GEN_80; // @[ICache.scala 57:28 ICache.scala 57:28]
  wire [52:0] _GEN_82 = 5'h12 == index_addr ? tag2_18 : _GEN_81; // @[ICache.scala 57:28 ICache.scala 57:28]
  wire [52:0] _GEN_83 = 5'h13 == index_addr ? tag2_19 : _GEN_82; // @[ICache.scala 57:28 ICache.scala 57:28]
  wire [52:0] _GEN_84 = 5'h14 == index_addr ? tag2_20 : _GEN_83; // @[ICache.scala 57:28 ICache.scala 57:28]
  wire [52:0] _GEN_85 = 5'h15 == index_addr ? tag2_21 : _GEN_84; // @[ICache.scala 57:28 ICache.scala 57:28]
  wire [52:0] _GEN_86 = 5'h16 == index_addr ? tag2_22 : _GEN_85; // @[ICache.scala 57:28 ICache.scala 57:28]
  wire [52:0] _GEN_87 = 5'h17 == index_addr ? tag2_23 : _GEN_86; // @[ICache.scala 57:28 ICache.scala 57:28]
  wire [52:0] _GEN_88 = 5'h18 == index_addr ? tag2_24 : _GEN_87; // @[ICache.scala 57:28 ICache.scala 57:28]
  wire [52:0] _GEN_89 = 5'h19 == index_addr ? tag2_25 : _GEN_88; // @[ICache.scala 57:28 ICache.scala 57:28]
  wire [52:0] _GEN_90 = 5'h1a == index_addr ? tag2_26 : _GEN_89; // @[ICache.scala 57:28 ICache.scala 57:28]
  wire [52:0] _GEN_91 = 5'h1b == index_addr ? tag2_27 : _GEN_90; // @[ICache.scala 57:28 ICache.scala 57:28]
  wire [52:0] _GEN_92 = 5'h1c == index_addr ? tag2_28 : _GEN_91; // @[ICache.scala 57:28 ICache.scala 57:28]
  wire [52:0] _GEN_93 = 5'h1d == index_addr ? tag2_29 : _GEN_92; // @[ICache.scala 57:28 ICache.scala 57:28]
  wire [52:0] _GEN_94 = 5'h1e == index_addr ? tag2_30 : _GEN_93; // @[ICache.scala 57:28 ICache.scala 57:28]
  wire [52:0] _GEN_95 = 5'h1f == index_addr ? tag2_31 : _GEN_94; // @[ICache.scala 57:28 ICache.scala 57:28]
  wire  _GEN_97 = 5'h1 == index_addr ? v2_1 : v2_0; // @[ICache.scala 57:67 ICache.scala 57:67]
  wire  _GEN_98 = 5'h2 == index_addr ? v2_2 : _GEN_97; // @[ICache.scala 57:67 ICache.scala 57:67]
  wire  _GEN_99 = 5'h3 == index_addr ? v2_3 : _GEN_98; // @[ICache.scala 57:67 ICache.scala 57:67]
  wire  _GEN_100 = 5'h4 == index_addr ? v2_4 : _GEN_99; // @[ICache.scala 57:67 ICache.scala 57:67]
  wire  _GEN_101 = 5'h5 == index_addr ? v2_5 : _GEN_100; // @[ICache.scala 57:67 ICache.scala 57:67]
  wire  _GEN_102 = 5'h6 == index_addr ? v2_6 : _GEN_101; // @[ICache.scala 57:67 ICache.scala 57:67]
  wire  _GEN_103 = 5'h7 == index_addr ? v2_7 : _GEN_102; // @[ICache.scala 57:67 ICache.scala 57:67]
  wire  _GEN_104 = 5'h8 == index_addr ? v2_8 : _GEN_103; // @[ICache.scala 57:67 ICache.scala 57:67]
  wire  _GEN_105 = 5'h9 == index_addr ? v2_9 : _GEN_104; // @[ICache.scala 57:67 ICache.scala 57:67]
  wire  _GEN_106 = 5'ha == index_addr ? v2_10 : _GEN_105; // @[ICache.scala 57:67 ICache.scala 57:67]
  wire  _GEN_107 = 5'hb == index_addr ? v2_11 : _GEN_106; // @[ICache.scala 57:67 ICache.scala 57:67]
  wire  _GEN_108 = 5'hc == index_addr ? v2_12 : _GEN_107; // @[ICache.scala 57:67 ICache.scala 57:67]
  wire  _GEN_109 = 5'hd == index_addr ? v2_13 : _GEN_108; // @[ICache.scala 57:67 ICache.scala 57:67]
  wire  _GEN_110 = 5'he == index_addr ? v2_14 : _GEN_109; // @[ICache.scala 57:67 ICache.scala 57:67]
  wire  _GEN_111 = 5'hf == index_addr ? v2_15 : _GEN_110; // @[ICache.scala 57:67 ICache.scala 57:67]
  wire  _GEN_112 = 5'h10 == index_addr ? v2_16 : _GEN_111; // @[ICache.scala 57:67 ICache.scala 57:67]
  wire  _GEN_113 = 5'h11 == index_addr ? v2_17 : _GEN_112; // @[ICache.scala 57:67 ICache.scala 57:67]
  wire  _GEN_114 = 5'h12 == index_addr ? v2_18 : _GEN_113; // @[ICache.scala 57:67 ICache.scala 57:67]
  wire  _GEN_115 = 5'h13 == index_addr ? v2_19 : _GEN_114; // @[ICache.scala 57:67 ICache.scala 57:67]
  wire  _GEN_116 = 5'h14 == index_addr ? v2_20 : _GEN_115; // @[ICache.scala 57:67 ICache.scala 57:67]
  wire  _GEN_117 = 5'h15 == index_addr ? v2_21 : _GEN_116; // @[ICache.scala 57:67 ICache.scala 57:67]
  wire  _GEN_118 = 5'h16 == index_addr ? v2_22 : _GEN_117; // @[ICache.scala 57:67 ICache.scala 57:67]
  wire  _GEN_119 = 5'h17 == index_addr ? v2_23 : _GEN_118; // @[ICache.scala 57:67 ICache.scala 57:67]
  wire  _GEN_120 = 5'h18 == index_addr ? v2_24 : _GEN_119; // @[ICache.scala 57:67 ICache.scala 57:67]
  wire  _GEN_121 = 5'h19 == index_addr ? v2_25 : _GEN_120; // @[ICache.scala 57:67 ICache.scala 57:67]
  wire  _GEN_122 = 5'h1a == index_addr ? v2_26 : _GEN_121; // @[ICache.scala 57:67 ICache.scala 57:67]
  wire  _GEN_123 = 5'h1b == index_addr ? v2_27 : _GEN_122; // @[ICache.scala 57:67 ICache.scala 57:67]
  wire  _GEN_124 = 5'h1c == index_addr ? v2_28 : _GEN_123; // @[ICache.scala 57:67 ICache.scala 57:67]
  wire  _GEN_125 = 5'h1d == index_addr ? v2_29 : _GEN_124; // @[ICache.scala 57:67 ICache.scala 57:67]
  wire  _GEN_126 = 5'h1e == index_addr ? v2_30 : _GEN_125; // @[ICache.scala 57:67 ICache.scala 57:67]
  wire  _GEN_127 = 5'h1f == index_addr ? v2_31 : _GEN_126; // @[ICache.scala 57:67 ICache.scala 57:67]
  wire  hit2 = tag_addr == _GEN_95 & _GEN_127; // @[ICache.scala 57:49]
  wire [8:0] _data1_T = {offset_addr, 3'h0}; // @[ICache.scala 58:55]
  wire [511:0] _GEN_129 = 5'h1 == index_addr ? block1_1 : block1_0; // @[ICache.scala 58:39 ICache.scala 58:39]
  wire [511:0] _GEN_130 = 5'h2 == index_addr ? block1_2 : _GEN_129; // @[ICache.scala 58:39 ICache.scala 58:39]
  wire [511:0] _GEN_131 = 5'h3 == index_addr ? block1_3 : _GEN_130; // @[ICache.scala 58:39 ICache.scala 58:39]
  wire [511:0] _GEN_132 = 5'h4 == index_addr ? block1_4 : _GEN_131; // @[ICache.scala 58:39 ICache.scala 58:39]
  wire [511:0] _GEN_133 = 5'h5 == index_addr ? block1_5 : _GEN_132; // @[ICache.scala 58:39 ICache.scala 58:39]
  wire [511:0] _GEN_134 = 5'h6 == index_addr ? block1_6 : _GEN_133; // @[ICache.scala 58:39 ICache.scala 58:39]
  wire [511:0] _GEN_135 = 5'h7 == index_addr ? block1_7 : _GEN_134; // @[ICache.scala 58:39 ICache.scala 58:39]
  wire [511:0] _GEN_136 = 5'h8 == index_addr ? block1_8 : _GEN_135; // @[ICache.scala 58:39 ICache.scala 58:39]
  wire [511:0] _GEN_137 = 5'h9 == index_addr ? block1_9 : _GEN_136; // @[ICache.scala 58:39 ICache.scala 58:39]
  wire [511:0] _GEN_138 = 5'ha == index_addr ? block1_10 : _GEN_137; // @[ICache.scala 58:39 ICache.scala 58:39]
  wire [511:0] _GEN_139 = 5'hb == index_addr ? block1_11 : _GEN_138; // @[ICache.scala 58:39 ICache.scala 58:39]
  wire [511:0] _GEN_140 = 5'hc == index_addr ? block1_12 : _GEN_139; // @[ICache.scala 58:39 ICache.scala 58:39]
  wire [511:0] _GEN_141 = 5'hd == index_addr ? block1_13 : _GEN_140; // @[ICache.scala 58:39 ICache.scala 58:39]
  wire [511:0] _GEN_142 = 5'he == index_addr ? block1_14 : _GEN_141; // @[ICache.scala 58:39 ICache.scala 58:39]
  wire [511:0] _GEN_143 = 5'hf == index_addr ? block1_15 : _GEN_142; // @[ICache.scala 58:39 ICache.scala 58:39]
  wire [511:0] _GEN_144 = 5'h10 == index_addr ? block1_16 : _GEN_143; // @[ICache.scala 58:39 ICache.scala 58:39]
  wire [511:0] _GEN_145 = 5'h11 == index_addr ? block1_17 : _GEN_144; // @[ICache.scala 58:39 ICache.scala 58:39]
  wire [511:0] _GEN_146 = 5'h12 == index_addr ? block1_18 : _GEN_145; // @[ICache.scala 58:39 ICache.scala 58:39]
  wire [511:0] _GEN_147 = 5'h13 == index_addr ? block1_19 : _GEN_146; // @[ICache.scala 58:39 ICache.scala 58:39]
  wire [511:0] _GEN_148 = 5'h14 == index_addr ? block1_20 : _GEN_147; // @[ICache.scala 58:39 ICache.scala 58:39]
  wire [511:0] _GEN_149 = 5'h15 == index_addr ? block1_21 : _GEN_148; // @[ICache.scala 58:39 ICache.scala 58:39]
  wire [511:0] _GEN_150 = 5'h16 == index_addr ? block1_22 : _GEN_149; // @[ICache.scala 58:39 ICache.scala 58:39]
  wire [511:0] _GEN_151 = 5'h17 == index_addr ? block1_23 : _GEN_150; // @[ICache.scala 58:39 ICache.scala 58:39]
  wire [511:0] _GEN_152 = 5'h18 == index_addr ? block1_24 : _GEN_151; // @[ICache.scala 58:39 ICache.scala 58:39]
  wire [511:0] _GEN_153 = 5'h19 == index_addr ? block1_25 : _GEN_152; // @[ICache.scala 58:39 ICache.scala 58:39]
  wire [511:0] _GEN_154 = 5'h1a == index_addr ? block1_26 : _GEN_153; // @[ICache.scala 58:39 ICache.scala 58:39]
  wire [511:0] _GEN_155 = 5'h1b == index_addr ? block1_27 : _GEN_154; // @[ICache.scala 58:39 ICache.scala 58:39]
  wire [511:0] _GEN_156 = 5'h1c == index_addr ? block1_28 : _GEN_155; // @[ICache.scala 58:39 ICache.scala 58:39]
  wire [511:0] _GEN_157 = 5'h1d == index_addr ? block1_29 : _GEN_156; // @[ICache.scala 58:39 ICache.scala 58:39]
  wire [511:0] _GEN_158 = 5'h1e == index_addr ? block1_30 : _GEN_157; // @[ICache.scala 58:39 ICache.scala 58:39]
  wire [511:0] _GEN_159 = 5'h1f == index_addr ? block1_31 : _GEN_158; // @[ICache.scala 58:39 ICache.scala 58:39]
  wire [511:0] _data1_T_1 = _GEN_159 >> _data1_T; // @[ICache.scala 58:39]
  wire [31:0] data1 = _data1_T_1[31:0]; // @[ICache.scala 58:61]
  wire [511:0] _GEN_161 = 5'h1 == index_addr ? block2_1 : block2_0; // @[ICache.scala 59:39 ICache.scala 59:39]
  wire [511:0] _GEN_162 = 5'h2 == index_addr ? block2_2 : _GEN_161; // @[ICache.scala 59:39 ICache.scala 59:39]
  wire [511:0] _GEN_163 = 5'h3 == index_addr ? block2_3 : _GEN_162; // @[ICache.scala 59:39 ICache.scala 59:39]
  wire [511:0] _GEN_164 = 5'h4 == index_addr ? block2_4 : _GEN_163; // @[ICache.scala 59:39 ICache.scala 59:39]
  wire [511:0] _GEN_165 = 5'h5 == index_addr ? block2_5 : _GEN_164; // @[ICache.scala 59:39 ICache.scala 59:39]
  wire [511:0] _GEN_166 = 5'h6 == index_addr ? block2_6 : _GEN_165; // @[ICache.scala 59:39 ICache.scala 59:39]
  wire [511:0] _GEN_167 = 5'h7 == index_addr ? block2_7 : _GEN_166; // @[ICache.scala 59:39 ICache.scala 59:39]
  wire [511:0] _GEN_168 = 5'h8 == index_addr ? block2_8 : _GEN_167; // @[ICache.scala 59:39 ICache.scala 59:39]
  wire [511:0] _GEN_169 = 5'h9 == index_addr ? block2_9 : _GEN_168; // @[ICache.scala 59:39 ICache.scala 59:39]
  wire [511:0] _GEN_170 = 5'ha == index_addr ? block2_10 : _GEN_169; // @[ICache.scala 59:39 ICache.scala 59:39]
  wire [511:0] _GEN_171 = 5'hb == index_addr ? block2_11 : _GEN_170; // @[ICache.scala 59:39 ICache.scala 59:39]
  wire [511:0] _GEN_172 = 5'hc == index_addr ? block2_12 : _GEN_171; // @[ICache.scala 59:39 ICache.scala 59:39]
  wire [511:0] _GEN_173 = 5'hd == index_addr ? block2_13 : _GEN_172; // @[ICache.scala 59:39 ICache.scala 59:39]
  wire [511:0] _GEN_174 = 5'he == index_addr ? block2_14 : _GEN_173; // @[ICache.scala 59:39 ICache.scala 59:39]
  wire [511:0] _GEN_175 = 5'hf == index_addr ? block2_15 : _GEN_174; // @[ICache.scala 59:39 ICache.scala 59:39]
  wire [511:0] _GEN_176 = 5'h10 == index_addr ? block2_16 : _GEN_175; // @[ICache.scala 59:39 ICache.scala 59:39]
  wire [511:0] _GEN_177 = 5'h11 == index_addr ? block2_17 : _GEN_176; // @[ICache.scala 59:39 ICache.scala 59:39]
  wire [511:0] _GEN_178 = 5'h12 == index_addr ? block2_18 : _GEN_177; // @[ICache.scala 59:39 ICache.scala 59:39]
  wire [511:0] _GEN_179 = 5'h13 == index_addr ? block2_19 : _GEN_178; // @[ICache.scala 59:39 ICache.scala 59:39]
  wire [511:0] _GEN_180 = 5'h14 == index_addr ? block2_20 : _GEN_179; // @[ICache.scala 59:39 ICache.scala 59:39]
  wire [511:0] _GEN_181 = 5'h15 == index_addr ? block2_21 : _GEN_180; // @[ICache.scala 59:39 ICache.scala 59:39]
  wire [511:0] _GEN_182 = 5'h16 == index_addr ? block2_22 : _GEN_181; // @[ICache.scala 59:39 ICache.scala 59:39]
  wire [511:0] _GEN_183 = 5'h17 == index_addr ? block2_23 : _GEN_182; // @[ICache.scala 59:39 ICache.scala 59:39]
  wire [511:0] _GEN_184 = 5'h18 == index_addr ? block2_24 : _GEN_183; // @[ICache.scala 59:39 ICache.scala 59:39]
  wire [511:0] _GEN_185 = 5'h19 == index_addr ? block2_25 : _GEN_184; // @[ICache.scala 59:39 ICache.scala 59:39]
  wire [511:0] _GEN_186 = 5'h1a == index_addr ? block2_26 : _GEN_185; // @[ICache.scala 59:39 ICache.scala 59:39]
  wire [511:0] _GEN_187 = 5'h1b == index_addr ? block2_27 : _GEN_186; // @[ICache.scala 59:39 ICache.scala 59:39]
  wire [511:0] _GEN_188 = 5'h1c == index_addr ? block2_28 : _GEN_187; // @[ICache.scala 59:39 ICache.scala 59:39]
  wire [511:0] _GEN_189 = 5'h1d == index_addr ? block2_29 : _GEN_188; // @[ICache.scala 59:39 ICache.scala 59:39]
  wire [511:0] _GEN_190 = 5'h1e == index_addr ? block2_30 : _GEN_189; // @[ICache.scala 59:39 ICache.scala 59:39]
  wire [511:0] _GEN_191 = 5'h1f == index_addr ? block2_31 : _GEN_190; // @[ICache.scala 59:39 ICache.scala 59:39]
  wire [511:0] _data2_T_1 = _GEN_191 >> _data1_T; // @[ICache.scala 59:39]
  wire [31:0] data2 = _data2_T_1[31:0]; // @[ICache.scala 59:61]
  wire  hit = hit1 | hit2; // @[ICache.scala 61:24]
  wire  _age1_T = hit1 ^ hit2; // @[ICache.scala 66:49]
  wire  _GEN_193 = 5'h1 == index_addr ? age1_1 : age1_0; // @[ICache.scala 66:28 ICache.scala 66:28]
  wire  _GEN_194 = 5'h2 == index_addr ? age1_2 : _GEN_193; // @[ICache.scala 66:28 ICache.scala 66:28]
  wire  _GEN_195 = 5'h3 == index_addr ? age1_3 : _GEN_194; // @[ICache.scala 66:28 ICache.scala 66:28]
  wire  _GEN_196 = 5'h4 == index_addr ? age1_4 : _GEN_195; // @[ICache.scala 66:28 ICache.scala 66:28]
  wire  _GEN_197 = 5'h5 == index_addr ? age1_5 : _GEN_196; // @[ICache.scala 66:28 ICache.scala 66:28]
  wire  _GEN_198 = 5'h6 == index_addr ? age1_6 : _GEN_197; // @[ICache.scala 66:28 ICache.scala 66:28]
  wire  _GEN_199 = 5'h7 == index_addr ? age1_7 : _GEN_198; // @[ICache.scala 66:28 ICache.scala 66:28]
  wire  _GEN_200 = 5'h8 == index_addr ? age1_8 : _GEN_199; // @[ICache.scala 66:28 ICache.scala 66:28]
  wire  _GEN_201 = 5'h9 == index_addr ? age1_9 : _GEN_200; // @[ICache.scala 66:28 ICache.scala 66:28]
  wire  _GEN_202 = 5'ha == index_addr ? age1_10 : _GEN_201; // @[ICache.scala 66:28 ICache.scala 66:28]
  wire  _GEN_203 = 5'hb == index_addr ? age1_11 : _GEN_202; // @[ICache.scala 66:28 ICache.scala 66:28]
  wire  _GEN_204 = 5'hc == index_addr ? age1_12 : _GEN_203; // @[ICache.scala 66:28 ICache.scala 66:28]
  wire  _GEN_205 = 5'hd == index_addr ? age1_13 : _GEN_204; // @[ICache.scala 66:28 ICache.scala 66:28]
  wire  _GEN_206 = 5'he == index_addr ? age1_14 : _GEN_205; // @[ICache.scala 66:28 ICache.scala 66:28]
  wire  _GEN_207 = 5'hf == index_addr ? age1_15 : _GEN_206; // @[ICache.scala 66:28 ICache.scala 66:28]
  wire  _GEN_208 = 5'h10 == index_addr ? age1_16 : _GEN_207; // @[ICache.scala 66:28 ICache.scala 66:28]
  wire  _GEN_209 = 5'h11 == index_addr ? age1_17 : _GEN_208; // @[ICache.scala 66:28 ICache.scala 66:28]
  wire  _GEN_210 = 5'h12 == index_addr ? age1_18 : _GEN_209; // @[ICache.scala 66:28 ICache.scala 66:28]
  wire  _GEN_211 = 5'h13 == index_addr ? age1_19 : _GEN_210; // @[ICache.scala 66:28 ICache.scala 66:28]
  wire  _GEN_212 = 5'h14 == index_addr ? age1_20 : _GEN_211; // @[ICache.scala 66:28 ICache.scala 66:28]
  wire  _GEN_213 = 5'h15 == index_addr ? age1_21 : _GEN_212; // @[ICache.scala 66:28 ICache.scala 66:28]
  wire  _GEN_214 = 5'h16 == index_addr ? age1_22 : _GEN_213; // @[ICache.scala 66:28 ICache.scala 66:28]
  wire  _GEN_215 = 5'h17 == index_addr ? age1_23 : _GEN_214; // @[ICache.scala 66:28 ICache.scala 66:28]
  wire  _GEN_216 = 5'h18 == index_addr ? age1_24 : _GEN_215; // @[ICache.scala 66:28 ICache.scala 66:28]
  wire  _GEN_217 = 5'h19 == index_addr ? age1_25 : _GEN_216; // @[ICache.scala 66:28 ICache.scala 66:28]
  wire  _GEN_218 = 5'h1a == index_addr ? age1_26 : _GEN_217; // @[ICache.scala 66:28 ICache.scala 66:28]
  wire  _GEN_219 = 5'h1b == index_addr ? age1_27 : _GEN_218; // @[ICache.scala 66:28 ICache.scala 66:28]
  wire  _GEN_220 = 5'h1c == index_addr ? age1_28 : _GEN_219; // @[ICache.scala 66:28 ICache.scala 66:28]
  wire  _GEN_221 = 5'h1d == index_addr ? age1_29 : _GEN_220; // @[ICache.scala 66:28 ICache.scala 66:28]
  wire  _GEN_222 = 5'h1e == index_addr ? age1_30 : _GEN_221; // @[ICache.scala 66:28 ICache.scala 66:28]
  wire  _GEN_223 = 5'h1f == index_addr ? age1_31 : _GEN_222; // @[ICache.scala 66:28 ICache.scala 66:28]
  wire  _GEN_257 = 5'h1 == index_addr ? age2_1 : age2_0; // @[ICache.scala 67:28 ICache.scala 67:28]
  wire  _GEN_258 = 5'h2 == index_addr ? age2_2 : _GEN_257; // @[ICache.scala 67:28 ICache.scala 67:28]
  wire  _GEN_259 = 5'h3 == index_addr ? age2_3 : _GEN_258; // @[ICache.scala 67:28 ICache.scala 67:28]
  wire  _GEN_260 = 5'h4 == index_addr ? age2_4 : _GEN_259; // @[ICache.scala 67:28 ICache.scala 67:28]
  wire  _GEN_261 = 5'h5 == index_addr ? age2_5 : _GEN_260; // @[ICache.scala 67:28 ICache.scala 67:28]
  wire  _GEN_262 = 5'h6 == index_addr ? age2_6 : _GEN_261; // @[ICache.scala 67:28 ICache.scala 67:28]
  wire  _GEN_263 = 5'h7 == index_addr ? age2_7 : _GEN_262; // @[ICache.scala 67:28 ICache.scala 67:28]
  wire  _GEN_264 = 5'h8 == index_addr ? age2_8 : _GEN_263; // @[ICache.scala 67:28 ICache.scala 67:28]
  wire  _GEN_265 = 5'h9 == index_addr ? age2_9 : _GEN_264; // @[ICache.scala 67:28 ICache.scala 67:28]
  wire  _GEN_266 = 5'ha == index_addr ? age2_10 : _GEN_265; // @[ICache.scala 67:28 ICache.scala 67:28]
  wire  _GEN_267 = 5'hb == index_addr ? age2_11 : _GEN_266; // @[ICache.scala 67:28 ICache.scala 67:28]
  wire  _GEN_268 = 5'hc == index_addr ? age2_12 : _GEN_267; // @[ICache.scala 67:28 ICache.scala 67:28]
  wire  _GEN_269 = 5'hd == index_addr ? age2_13 : _GEN_268; // @[ICache.scala 67:28 ICache.scala 67:28]
  wire  _GEN_270 = 5'he == index_addr ? age2_14 : _GEN_269; // @[ICache.scala 67:28 ICache.scala 67:28]
  wire  _GEN_271 = 5'hf == index_addr ? age2_15 : _GEN_270; // @[ICache.scala 67:28 ICache.scala 67:28]
  wire  _GEN_272 = 5'h10 == index_addr ? age2_16 : _GEN_271; // @[ICache.scala 67:28 ICache.scala 67:28]
  wire  _GEN_273 = 5'h11 == index_addr ? age2_17 : _GEN_272; // @[ICache.scala 67:28 ICache.scala 67:28]
  wire  _GEN_274 = 5'h12 == index_addr ? age2_18 : _GEN_273; // @[ICache.scala 67:28 ICache.scala 67:28]
  wire  _GEN_275 = 5'h13 == index_addr ? age2_19 : _GEN_274; // @[ICache.scala 67:28 ICache.scala 67:28]
  wire  _GEN_276 = 5'h14 == index_addr ? age2_20 : _GEN_275; // @[ICache.scala 67:28 ICache.scala 67:28]
  wire  _GEN_277 = 5'h15 == index_addr ? age2_21 : _GEN_276; // @[ICache.scala 67:28 ICache.scala 67:28]
  wire  _GEN_278 = 5'h16 == index_addr ? age2_22 : _GEN_277; // @[ICache.scala 67:28 ICache.scala 67:28]
  wire  _GEN_279 = 5'h17 == index_addr ? age2_23 : _GEN_278; // @[ICache.scala 67:28 ICache.scala 67:28]
  wire  _GEN_280 = 5'h18 == index_addr ? age2_24 : _GEN_279; // @[ICache.scala 67:28 ICache.scala 67:28]
  wire  _GEN_281 = 5'h19 == index_addr ? age2_25 : _GEN_280; // @[ICache.scala 67:28 ICache.scala 67:28]
  wire  _GEN_282 = 5'h1a == index_addr ? age2_26 : _GEN_281; // @[ICache.scala 67:28 ICache.scala 67:28]
  wire  _GEN_283 = 5'h1b == index_addr ? age2_27 : _GEN_282; // @[ICache.scala 67:28 ICache.scala 67:28]
  wire  _GEN_284 = 5'h1c == index_addr ? age2_28 : _GEN_283; // @[ICache.scala 67:28 ICache.scala 67:28]
  wire  _GEN_285 = 5'h1d == index_addr ? age2_29 : _GEN_284; // @[ICache.scala 67:28 ICache.scala 67:28]
  wire  _GEN_286 = 5'h1e == index_addr ? age2_30 : _GEN_285; // @[ICache.scala 67:28 ICache.scala 67:28]
  wire  _GEN_287 = 5'h1f == index_addr ? age2_31 : _GEN_286; // @[ICache.scala 67:28 ICache.scala 67:28]
  reg [31:0] io_imem_data_REG; // @[ICache.scala 69:31]
  reg  io_imem_data_ok_REG; // @[ICache.scala 70:31]
  reg  state; // @[ICache.scala 75:24]
  wire  _T = ~state; // @[Conditional.scala 37:30]
  wire  _GEN_320 = ~hit | state; // @[ICache.scala 79:38 ICache.scala 79:45 ICache.scala 75:24]
  wire [1:0] age = {_GEN_287,_GEN_223}; // @[Cat.scala 30:58]
  wire  updateway2 = age == 2'h1; // @[ICache.scala 92:26]
  wire  updateway1 = ~updateway2; // @[ICache.scala 93:22]
  wire  update = state & io_axi_valid; // @[ICache.scala 94:33]
  wire  _block1_T = update & updateway1; // @[ICache.scala 95:40]
  wire  _block2_T = update & updateway2; // @[ICache.scala 98:40]
  assign io_imem_data = io_imem_data_REG; // @[ICache.scala 69:21]
  assign io_imem_data_ok = io_imem_data_ok_REG; // @[ICache.scala 70:21]
  assign io_axi_req = state; // @[ICache.scala 87:28]
  assign io_axi_addr = io_imem_addr & 64'hffffffffffffffc0; // @[ICache.scala 88:35]
  always @(posedge clock) begin
    if (reset) begin // @[ICache.scala 47:26]
      v1_0 <= 1'h0; // @[ICache.scala 47:26]
    end else if (5'h0 == index_addr) begin // @[ICache.scala 97:26]
      v1_0 <= _block1_T | _GEN_63; // @[ICache.scala 97:26]
    end
    if (reset) begin // @[ICache.scala 47:26]
      v1_1 <= 1'h0; // @[ICache.scala 47:26]
    end else if (5'h1 == index_addr) begin // @[ICache.scala 97:26]
      v1_1 <= _block1_T | _GEN_63; // @[ICache.scala 97:26]
    end
    if (reset) begin // @[ICache.scala 47:26]
      v1_2 <= 1'h0; // @[ICache.scala 47:26]
    end else if (5'h2 == index_addr) begin // @[ICache.scala 97:26]
      v1_2 <= _block1_T | _GEN_63; // @[ICache.scala 97:26]
    end
    if (reset) begin // @[ICache.scala 47:26]
      v1_3 <= 1'h0; // @[ICache.scala 47:26]
    end else if (5'h3 == index_addr) begin // @[ICache.scala 97:26]
      v1_3 <= _block1_T | _GEN_63; // @[ICache.scala 97:26]
    end
    if (reset) begin // @[ICache.scala 47:26]
      v1_4 <= 1'h0; // @[ICache.scala 47:26]
    end else if (5'h4 == index_addr) begin // @[ICache.scala 97:26]
      v1_4 <= _block1_T | _GEN_63; // @[ICache.scala 97:26]
    end
    if (reset) begin // @[ICache.scala 47:26]
      v1_5 <= 1'h0; // @[ICache.scala 47:26]
    end else if (5'h5 == index_addr) begin // @[ICache.scala 97:26]
      v1_5 <= _block1_T | _GEN_63; // @[ICache.scala 97:26]
    end
    if (reset) begin // @[ICache.scala 47:26]
      v1_6 <= 1'h0; // @[ICache.scala 47:26]
    end else if (5'h6 == index_addr) begin // @[ICache.scala 97:26]
      v1_6 <= _block1_T | _GEN_63; // @[ICache.scala 97:26]
    end
    if (reset) begin // @[ICache.scala 47:26]
      v1_7 <= 1'h0; // @[ICache.scala 47:26]
    end else if (5'h7 == index_addr) begin // @[ICache.scala 97:26]
      v1_7 <= _block1_T | _GEN_63; // @[ICache.scala 97:26]
    end
    if (reset) begin // @[ICache.scala 47:26]
      v1_8 <= 1'h0; // @[ICache.scala 47:26]
    end else if (5'h8 == index_addr) begin // @[ICache.scala 97:26]
      v1_8 <= _block1_T | _GEN_63; // @[ICache.scala 97:26]
    end
    if (reset) begin // @[ICache.scala 47:26]
      v1_9 <= 1'h0; // @[ICache.scala 47:26]
    end else if (5'h9 == index_addr) begin // @[ICache.scala 97:26]
      v1_9 <= _block1_T | _GEN_63; // @[ICache.scala 97:26]
    end
    if (reset) begin // @[ICache.scala 47:26]
      v1_10 <= 1'h0; // @[ICache.scala 47:26]
    end else if (5'ha == index_addr) begin // @[ICache.scala 97:26]
      v1_10 <= _block1_T | _GEN_63; // @[ICache.scala 97:26]
    end
    if (reset) begin // @[ICache.scala 47:26]
      v1_11 <= 1'h0; // @[ICache.scala 47:26]
    end else if (5'hb == index_addr) begin // @[ICache.scala 97:26]
      v1_11 <= _block1_T | _GEN_63; // @[ICache.scala 97:26]
    end
    if (reset) begin // @[ICache.scala 47:26]
      v1_12 <= 1'h0; // @[ICache.scala 47:26]
    end else if (5'hc == index_addr) begin // @[ICache.scala 97:26]
      v1_12 <= _block1_T | _GEN_63; // @[ICache.scala 97:26]
    end
    if (reset) begin // @[ICache.scala 47:26]
      v1_13 <= 1'h0; // @[ICache.scala 47:26]
    end else if (5'hd == index_addr) begin // @[ICache.scala 97:26]
      v1_13 <= _block1_T | _GEN_63; // @[ICache.scala 97:26]
    end
    if (reset) begin // @[ICache.scala 47:26]
      v1_14 <= 1'h0; // @[ICache.scala 47:26]
    end else if (5'he == index_addr) begin // @[ICache.scala 97:26]
      v1_14 <= _block1_T | _GEN_63; // @[ICache.scala 97:26]
    end
    if (reset) begin // @[ICache.scala 47:26]
      v1_15 <= 1'h0; // @[ICache.scala 47:26]
    end else if (5'hf == index_addr) begin // @[ICache.scala 97:26]
      v1_15 <= _block1_T | _GEN_63; // @[ICache.scala 97:26]
    end
    if (reset) begin // @[ICache.scala 47:26]
      v1_16 <= 1'h0; // @[ICache.scala 47:26]
    end else if (5'h10 == index_addr) begin // @[ICache.scala 97:26]
      v1_16 <= _block1_T | _GEN_63; // @[ICache.scala 97:26]
    end
    if (reset) begin // @[ICache.scala 47:26]
      v1_17 <= 1'h0; // @[ICache.scala 47:26]
    end else if (5'h11 == index_addr) begin // @[ICache.scala 97:26]
      v1_17 <= _block1_T | _GEN_63; // @[ICache.scala 97:26]
    end
    if (reset) begin // @[ICache.scala 47:26]
      v1_18 <= 1'h0; // @[ICache.scala 47:26]
    end else if (5'h12 == index_addr) begin // @[ICache.scala 97:26]
      v1_18 <= _block1_T | _GEN_63; // @[ICache.scala 97:26]
    end
    if (reset) begin // @[ICache.scala 47:26]
      v1_19 <= 1'h0; // @[ICache.scala 47:26]
    end else if (5'h13 == index_addr) begin // @[ICache.scala 97:26]
      v1_19 <= _block1_T | _GEN_63; // @[ICache.scala 97:26]
    end
    if (reset) begin // @[ICache.scala 47:26]
      v1_20 <= 1'h0; // @[ICache.scala 47:26]
    end else if (5'h14 == index_addr) begin // @[ICache.scala 97:26]
      v1_20 <= _block1_T | _GEN_63; // @[ICache.scala 97:26]
    end
    if (reset) begin // @[ICache.scala 47:26]
      v1_21 <= 1'h0; // @[ICache.scala 47:26]
    end else if (5'h15 == index_addr) begin // @[ICache.scala 97:26]
      v1_21 <= _block1_T | _GEN_63; // @[ICache.scala 97:26]
    end
    if (reset) begin // @[ICache.scala 47:26]
      v1_22 <= 1'h0; // @[ICache.scala 47:26]
    end else if (5'h16 == index_addr) begin // @[ICache.scala 97:26]
      v1_22 <= _block1_T | _GEN_63; // @[ICache.scala 97:26]
    end
    if (reset) begin // @[ICache.scala 47:26]
      v1_23 <= 1'h0; // @[ICache.scala 47:26]
    end else if (5'h17 == index_addr) begin // @[ICache.scala 97:26]
      v1_23 <= _block1_T | _GEN_63; // @[ICache.scala 97:26]
    end
    if (reset) begin // @[ICache.scala 47:26]
      v1_24 <= 1'h0; // @[ICache.scala 47:26]
    end else if (5'h18 == index_addr) begin // @[ICache.scala 97:26]
      v1_24 <= _block1_T | _GEN_63; // @[ICache.scala 97:26]
    end
    if (reset) begin // @[ICache.scala 47:26]
      v1_25 <= 1'h0; // @[ICache.scala 47:26]
    end else if (5'h19 == index_addr) begin // @[ICache.scala 97:26]
      v1_25 <= _block1_T | _GEN_63; // @[ICache.scala 97:26]
    end
    if (reset) begin // @[ICache.scala 47:26]
      v1_26 <= 1'h0; // @[ICache.scala 47:26]
    end else if (5'h1a == index_addr) begin // @[ICache.scala 97:26]
      v1_26 <= _block1_T | _GEN_63; // @[ICache.scala 97:26]
    end
    if (reset) begin // @[ICache.scala 47:26]
      v1_27 <= 1'h0; // @[ICache.scala 47:26]
    end else if (5'h1b == index_addr) begin // @[ICache.scala 97:26]
      v1_27 <= _block1_T | _GEN_63; // @[ICache.scala 97:26]
    end
    if (reset) begin // @[ICache.scala 47:26]
      v1_28 <= 1'h0; // @[ICache.scala 47:26]
    end else if (5'h1c == index_addr) begin // @[ICache.scala 97:26]
      v1_28 <= _block1_T | _GEN_63; // @[ICache.scala 97:26]
    end
    if (reset) begin // @[ICache.scala 47:26]
      v1_29 <= 1'h0; // @[ICache.scala 47:26]
    end else if (5'h1d == index_addr) begin // @[ICache.scala 97:26]
      v1_29 <= _block1_T | _GEN_63; // @[ICache.scala 97:26]
    end
    if (reset) begin // @[ICache.scala 47:26]
      v1_30 <= 1'h0; // @[ICache.scala 47:26]
    end else if (5'h1e == index_addr) begin // @[ICache.scala 97:26]
      v1_30 <= _block1_T | _GEN_63; // @[ICache.scala 97:26]
    end
    if (reset) begin // @[ICache.scala 47:26]
      v1_31 <= 1'h0; // @[ICache.scala 47:26]
    end else if (5'h1f == index_addr) begin // @[ICache.scala 97:26]
      v1_31 <= _block1_T | _GEN_63; // @[ICache.scala 97:26]
    end
    if (reset) begin // @[ICache.scala 48:26]
      age1_0 <= 1'h0; // @[ICache.scala 48:26]
    end else if (5'h0 == index_addr) begin // @[ICache.scala 66:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 66:28]
        age1_0 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 66:28]
        age1_0 <= age1_31; // @[ICache.scala 66:28]
      end else begin
        age1_0 <= _GEN_222;
      end
    end
    if (reset) begin // @[ICache.scala 48:26]
      age1_1 <= 1'h0; // @[ICache.scala 48:26]
    end else if (5'h1 == index_addr) begin // @[ICache.scala 66:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 66:28]
        age1_1 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 66:28]
        age1_1 <= age1_31; // @[ICache.scala 66:28]
      end else begin
        age1_1 <= _GEN_222;
      end
    end
    if (reset) begin // @[ICache.scala 48:26]
      age1_2 <= 1'h0; // @[ICache.scala 48:26]
    end else if (5'h2 == index_addr) begin // @[ICache.scala 66:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 66:28]
        age1_2 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 66:28]
        age1_2 <= age1_31; // @[ICache.scala 66:28]
      end else begin
        age1_2 <= _GEN_222;
      end
    end
    if (reset) begin // @[ICache.scala 48:26]
      age1_3 <= 1'h0; // @[ICache.scala 48:26]
    end else if (5'h3 == index_addr) begin // @[ICache.scala 66:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 66:28]
        age1_3 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 66:28]
        age1_3 <= age1_31; // @[ICache.scala 66:28]
      end else begin
        age1_3 <= _GEN_222;
      end
    end
    if (reset) begin // @[ICache.scala 48:26]
      age1_4 <= 1'h0; // @[ICache.scala 48:26]
    end else if (5'h4 == index_addr) begin // @[ICache.scala 66:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 66:28]
        age1_4 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 66:28]
        age1_4 <= age1_31; // @[ICache.scala 66:28]
      end else begin
        age1_4 <= _GEN_222;
      end
    end
    if (reset) begin // @[ICache.scala 48:26]
      age1_5 <= 1'h0; // @[ICache.scala 48:26]
    end else if (5'h5 == index_addr) begin // @[ICache.scala 66:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 66:28]
        age1_5 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 66:28]
        age1_5 <= age1_31; // @[ICache.scala 66:28]
      end else begin
        age1_5 <= _GEN_222;
      end
    end
    if (reset) begin // @[ICache.scala 48:26]
      age1_6 <= 1'h0; // @[ICache.scala 48:26]
    end else if (5'h6 == index_addr) begin // @[ICache.scala 66:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 66:28]
        age1_6 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 66:28]
        age1_6 <= age1_31; // @[ICache.scala 66:28]
      end else begin
        age1_6 <= _GEN_222;
      end
    end
    if (reset) begin // @[ICache.scala 48:26]
      age1_7 <= 1'h0; // @[ICache.scala 48:26]
    end else if (5'h7 == index_addr) begin // @[ICache.scala 66:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 66:28]
        age1_7 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 66:28]
        age1_7 <= age1_31; // @[ICache.scala 66:28]
      end else begin
        age1_7 <= _GEN_222;
      end
    end
    if (reset) begin // @[ICache.scala 48:26]
      age1_8 <= 1'h0; // @[ICache.scala 48:26]
    end else if (5'h8 == index_addr) begin // @[ICache.scala 66:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 66:28]
        age1_8 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 66:28]
        age1_8 <= age1_31; // @[ICache.scala 66:28]
      end else begin
        age1_8 <= _GEN_222;
      end
    end
    if (reset) begin // @[ICache.scala 48:26]
      age1_9 <= 1'h0; // @[ICache.scala 48:26]
    end else if (5'h9 == index_addr) begin // @[ICache.scala 66:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 66:28]
        age1_9 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 66:28]
        age1_9 <= age1_31; // @[ICache.scala 66:28]
      end else begin
        age1_9 <= _GEN_222;
      end
    end
    if (reset) begin // @[ICache.scala 48:26]
      age1_10 <= 1'h0; // @[ICache.scala 48:26]
    end else if (5'ha == index_addr) begin // @[ICache.scala 66:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 66:28]
        age1_10 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 66:28]
        age1_10 <= age1_31; // @[ICache.scala 66:28]
      end else begin
        age1_10 <= _GEN_222;
      end
    end
    if (reset) begin // @[ICache.scala 48:26]
      age1_11 <= 1'h0; // @[ICache.scala 48:26]
    end else if (5'hb == index_addr) begin // @[ICache.scala 66:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 66:28]
        age1_11 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 66:28]
        age1_11 <= age1_31; // @[ICache.scala 66:28]
      end else begin
        age1_11 <= _GEN_222;
      end
    end
    if (reset) begin // @[ICache.scala 48:26]
      age1_12 <= 1'h0; // @[ICache.scala 48:26]
    end else if (5'hc == index_addr) begin // @[ICache.scala 66:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 66:28]
        age1_12 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 66:28]
        age1_12 <= age1_31; // @[ICache.scala 66:28]
      end else begin
        age1_12 <= _GEN_222;
      end
    end
    if (reset) begin // @[ICache.scala 48:26]
      age1_13 <= 1'h0; // @[ICache.scala 48:26]
    end else if (5'hd == index_addr) begin // @[ICache.scala 66:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 66:28]
        age1_13 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 66:28]
        age1_13 <= age1_31; // @[ICache.scala 66:28]
      end else begin
        age1_13 <= _GEN_222;
      end
    end
    if (reset) begin // @[ICache.scala 48:26]
      age1_14 <= 1'h0; // @[ICache.scala 48:26]
    end else if (5'he == index_addr) begin // @[ICache.scala 66:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 66:28]
        age1_14 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 66:28]
        age1_14 <= age1_31; // @[ICache.scala 66:28]
      end else begin
        age1_14 <= _GEN_222;
      end
    end
    if (reset) begin // @[ICache.scala 48:26]
      age1_15 <= 1'h0; // @[ICache.scala 48:26]
    end else if (5'hf == index_addr) begin // @[ICache.scala 66:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 66:28]
        age1_15 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 66:28]
        age1_15 <= age1_31; // @[ICache.scala 66:28]
      end else begin
        age1_15 <= _GEN_222;
      end
    end
    if (reset) begin // @[ICache.scala 48:26]
      age1_16 <= 1'h0; // @[ICache.scala 48:26]
    end else if (5'h10 == index_addr) begin // @[ICache.scala 66:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 66:28]
        age1_16 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 66:28]
        age1_16 <= age1_31; // @[ICache.scala 66:28]
      end else begin
        age1_16 <= _GEN_222;
      end
    end
    if (reset) begin // @[ICache.scala 48:26]
      age1_17 <= 1'h0; // @[ICache.scala 48:26]
    end else if (5'h11 == index_addr) begin // @[ICache.scala 66:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 66:28]
        age1_17 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 66:28]
        age1_17 <= age1_31; // @[ICache.scala 66:28]
      end else begin
        age1_17 <= _GEN_222;
      end
    end
    if (reset) begin // @[ICache.scala 48:26]
      age1_18 <= 1'h0; // @[ICache.scala 48:26]
    end else if (5'h12 == index_addr) begin // @[ICache.scala 66:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 66:28]
        age1_18 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 66:28]
        age1_18 <= age1_31; // @[ICache.scala 66:28]
      end else begin
        age1_18 <= _GEN_222;
      end
    end
    if (reset) begin // @[ICache.scala 48:26]
      age1_19 <= 1'h0; // @[ICache.scala 48:26]
    end else if (5'h13 == index_addr) begin // @[ICache.scala 66:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 66:28]
        age1_19 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 66:28]
        age1_19 <= age1_31; // @[ICache.scala 66:28]
      end else begin
        age1_19 <= _GEN_222;
      end
    end
    if (reset) begin // @[ICache.scala 48:26]
      age1_20 <= 1'h0; // @[ICache.scala 48:26]
    end else if (5'h14 == index_addr) begin // @[ICache.scala 66:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 66:28]
        age1_20 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 66:28]
        age1_20 <= age1_31; // @[ICache.scala 66:28]
      end else begin
        age1_20 <= _GEN_222;
      end
    end
    if (reset) begin // @[ICache.scala 48:26]
      age1_21 <= 1'h0; // @[ICache.scala 48:26]
    end else if (5'h15 == index_addr) begin // @[ICache.scala 66:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 66:28]
        age1_21 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 66:28]
        age1_21 <= age1_31; // @[ICache.scala 66:28]
      end else begin
        age1_21 <= _GEN_222;
      end
    end
    if (reset) begin // @[ICache.scala 48:26]
      age1_22 <= 1'h0; // @[ICache.scala 48:26]
    end else if (5'h16 == index_addr) begin // @[ICache.scala 66:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 66:28]
        age1_22 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 66:28]
        age1_22 <= age1_31; // @[ICache.scala 66:28]
      end else begin
        age1_22 <= _GEN_222;
      end
    end
    if (reset) begin // @[ICache.scala 48:26]
      age1_23 <= 1'h0; // @[ICache.scala 48:26]
    end else if (5'h17 == index_addr) begin // @[ICache.scala 66:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 66:28]
        age1_23 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 66:28]
        age1_23 <= age1_31; // @[ICache.scala 66:28]
      end else begin
        age1_23 <= _GEN_222;
      end
    end
    if (reset) begin // @[ICache.scala 48:26]
      age1_24 <= 1'h0; // @[ICache.scala 48:26]
    end else if (5'h18 == index_addr) begin // @[ICache.scala 66:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 66:28]
        age1_24 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 66:28]
        age1_24 <= age1_31; // @[ICache.scala 66:28]
      end else begin
        age1_24 <= _GEN_222;
      end
    end
    if (reset) begin // @[ICache.scala 48:26]
      age1_25 <= 1'h0; // @[ICache.scala 48:26]
    end else if (5'h19 == index_addr) begin // @[ICache.scala 66:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 66:28]
        age1_25 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 66:28]
        age1_25 <= age1_31; // @[ICache.scala 66:28]
      end else begin
        age1_25 <= _GEN_222;
      end
    end
    if (reset) begin // @[ICache.scala 48:26]
      age1_26 <= 1'h0; // @[ICache.scala 48:26]
    end else if (5'h1a == index_addr) begin // @[ICache.scala 66:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 66:28]
        age1_26 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 66:28]
        age1_26 <= age1_31; // @[ICache.scala 66:28]
      end else begin
        age1_26 <= _GEN_222;
      end
    end
    if (reset) begin // @[ICache.scala 48:26]
      age1_27 <= 1'h0; // @[ICache.scala 48:26]
    end else if (5'h1b == index_addr) begin // @[ICache.scala 66:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 66:28]
        age1_27 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 66:28]
        age1_27 <= age1_31; // @[ICache.scala 66:28]
      end else begin
        age1_27 <= _GEN_222;
      end
    end
    if (reset) begin // @[ICache.scala 48:26]
      age1_28 <= 1'h0; // @[ICache.scala 48:26]
    end else if (5'h1c == index_addr) begin // @[ICache.scala 66:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 66:28]
        age1_28 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 66:28]
        age1_28 <= age1_31; // @[ICache.scala 66:28]
      end else begin
        age1_28 <= _GEN_222;
      end
    end
    if (reset) begin // @[ICache.scala 48:26]
      age1_29 <= 1'h0; // @[ICache.scala 48:26]
    end else if (5'h1d == index_addr) begin // @[ICache.scala 66:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 66:28]
        age1_29 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 66:28]
        age1_29 <= age1_31; // @[ICache.scala 66:28]
      end else begin
        age1_29 <= _GEN_222;
      end
    end
    if (reset) begin // @[ICache.scala 48:26]
      age1_30 <= 1'h0; // @[ICache.scala 48:26]
    end else if (5'h1e == index_addr) begin // @[ICache.scala 66:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 66:28]
        age1_30 <= hit1;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 66:28]
        age1_30 <= age1_31; // @[ICache.scala 66:28]
      end else begin
        age1_30 <= _GEN_222;
      end
    end
    if (reset) begin // @[ICache.scala 48:26]
      age1_31 <= 1'h0; // @[ICache.scala 48:26]
    end else if (5'h1f == index_addr) begin // @[ICache.scala 66:22]
      if (hit1 ^ hit2) begin // @[ICache.scala 66:28]
        age1_31 <= hit1;
      end else if (!(5'h1f == index_addr)) begin // @[ICache.scala 66:28]
        age1_31 <= _GEN_222;
      end
    end
    if (reset) begin // @[ICache.scala 49:26]
      tag1_0 <= 53'h0; // @[ICache.scala 49:26]
    end else if (5'h0 == index_addr) begin // @[ICache.scala 96:26]
      if (_block1_T) begin // @[ICache.scala 96:32]
        tag1_0 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 56:28]
        tag1_0 <= tag1_31; // @[ICache.scala 56:28]
      end else begin
        tag1_0 <= _GEN_30;
      end
    end
    if (reset) begin // @[ICache.scala 49:26]
      tag1_1 <= 53'h0; // @[ICache.scala 49:26]
    end else if (5'h1 == index_addr) begin // @[ICache.scala 96:26]
      if (_block1_T) begin // @[ICache.scala 96:32]
        tag1_1 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 56:28]
        tag1_1 <= tag1_31; // @[ICache.scala 56:28]
      end else begin
        tag1_1 <= _GEN_30;
      end
    end
    if (reset) begin // @[ICache.scala 49:26]
      tag1_2 <= 53'h0; // @[ICache.scala 49:26]
    end else if (5'h2 == index_addr) begin // @[ICache.scala 96:26]
      if (_block1_T) begin // @[ICache.scala 96:32]
        tag1_2 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 56:28]
        tag1_2 <= tag1_31; // @[ICache.scala 56:28]
      end else begin
        tag1_2 <= _GEN_30;
      end
    end
    if (reset) begin // @[ICache.scala 49:26]
      tag1_3 <= 53'h0; // @[ICache.scala 49:26]
    end else if (5'h3 == index_addr) begin // @[ICache.scala 96:26]
      if (_block1_T) begin // @[ICache.scala 96:32]
        tag1_3 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 56:28]
        tag1_3 <= tag1_31; // @[ICache.scala 56:28]
      end else begin
        tag1_3 <= _GEN_30;
      end
    end
    if (reset) begin // @[ICache.scala 49:26]
      tag1_4 <= 53'h0; // @[ICache.scala 49:26]
    end else if (5'h4 == index_addr) begin // @[ICache.scala 96:26]
      if (_block1_T) begin // @[ICache.scala 96:32]
        tag1_4 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 56:28]
        tag1_4 <= tag1_31; // @[ICache.scala 56:28]
      end else begin
        tag1_4 <= _GEN_30;
      end
    end
    if (reset) begin // @[ICache.scala 49:26]
      tag1_5 <= 53'h0; // @[ICache.scala 49:26]
    end else if (5'h5 == index_addr) begin // @[ICache.scala 96:26]
      if (_block1_T) begin // @[ICache.scala 96:32]
        tag1_5 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 56:28]
        tag1_5 <= tag1_31; // @[ICache.scala 56:28]
      end else begin
        tag1_5 <= _GEN_30;
      end
    end
    if (reset) begin // @[ICache.scala 49:26]
      tag1_6 <= 53'h0; // @[ICache.scala 49:26]
    end else if (5'h6 == index_addr) begin // @[ICache.scala 96:26]
      if (_block1_T) begin // @[ICache.scala 96:32]
        tag1_6 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 56:28]
        tag1_6 <= tag1_31; // @[ICache.scala 56:28]
      end else begin
        tag1_6 <= _GEN_30;
      end
    end
    if (reset) begin // @[ICache.scala 49:26]
      tag1_7 <= 53'h0; // @[ICache.scala 49:26]
    end else if (5'h7 == index_addr) begin // @[ICache.scala 96:26]
      if (_block1_T) begin // @[ICache.scala 96:32]
        tag1_7 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 56:28]
        tag1_7 <= tag1_31; // @[ICache.scala 56:28]
      end else begin
        tag1_7 <= _GEN_30;
      end
    end
    if (reset) begin // @[ICache.scala 49:26]
      tag1_8 <= 53'h0; // @[ICache.scala 49:26]
    end else if (5'h8 == index_addr) begin // @[ICache.scala 96:26]
      if (_block1_T) begin // @[ICache.scala 96:32]
        tag1_8 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 56:28]
        tag1_8 <= tag1_31; // @[ICache.scala 56:28]
      end else begin
        tag1_8 <= _GEN_30;
      end
    end
    if (reset) begin // @[ICache.scala 49:26]
      tag1_9 <= 53'h0; // @[ICache.scala 49:26]
    end else if (5'h9 == index_addr) begin // @[ICache.scala 96:26]
      if (_block1_T) begin // @[ICache.scala 96:32]
        tag1_9 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 56:28]
        tag1_9 <= tag1_31; // @[ICache.scala 56:28]
      end else begin
        tag1_9 <= _GEN_30;
      end
    end
    if (reset) begin // @[ICache.scala 49:26]
      tag1_10 <= 53'h0; // @[ICache.scala 49:26]
    end else if (5'ha == index_addr) begin // @[ICache.scala 96:26]
      if (_block1_T) begin // @[ICache.scala 96:32]
        tag1_10 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 56:28]
        tag1_10 <= tag1_31; // @[ICache.scala 56:28]
      end else begin
        tag1_10 <= _GEN_30;
      end
    end
    if (reset) begin // @[ICache.scala 49:26]
      tag1_11 <= 53'h0; // @[ICache.scala 49:26]
    end else if (5'hb == index_addr) begin // @[ICache.scala 96:26]
      if (_block1_T) begin // @[ICache.scala 96:32]
        tag1_11 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 56:28]
        tag1_11 <= tag1_31; // @[ICache.scala 56:28]
      end else begin
        tag1_11 <= _GEN_30;
      end
    end
    if (reset) begin // @[ICache.scala 49:26]
      tag1_12 <= 53'h0; // @[ICache.scala 49:26]
    end else if (5'hc == index_addr) begin // @[ICache.scala 96:26]
      if (_block1_T) begin // @[ICache.scala 96:32]
        tag1_12 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 56:28]
        tag1_12 <= tag1_31; // @[ICache.scala 56:28]
      end else begin
        tag1_12 <= _GEN_30;
      end
    end
    if (reset) begin // @[ICache.scala 49:26]
      tag1_13 <= 53'h0; // @[ICache.scala 49:26]
    end else if (5'hd == index_addr) begin // @[ICache.scala 96:26]
      if (_block1_T) begin // @[ICache.scala 96:32]
        tag1_13 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 56:28]
        tag1_13 <= tag1_31; // @[ICache.scala 56:28]
      end else begin
        tag1_13 <= _GEN_30;
      end
    end
    if (reset) begin // @[ICache.scala 49:26]
      tag1_14 <= 53'h0; // @[ICache.scala 49:26]
    end else if (5'he == index_addr) begin // @[ICache.scala 96:26]
      if (_block1_T) begin // @[ICache.scala 96:32]
        tag1_14 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 56:28]
        tag1_14 <= tag1_31; // @[ICache.scala 56:28]
      end else begin
        tag1_14 <= _GEN_30;
      end
    end
    if (reset) begin // @[ICache.scala 49:26]
      tag1_15 <= 53'h0; // @[ICache.scala 49:26]
    end else if (5'hf == index_addr) begin // @[ICache.scala 96:26]
      if (_block1_T) begin // @[ICache.scala 96:32]
        tag1_15 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 56:28]
        tag1_15 <= tag1_31; // @[ICache.scala 56:28]
      end else begin
        tag1_15 <= _GEN_30;
      end
    end
    if (reset) begin // @[ICache.scala 49:26]
      tag1_16 <= 53'h0; // @[ICache.scala 49:26]
    end else if (5'h10 == index_addr) begin // @[ICache.scala 96:26]
      if (_block1_T) begin // @[ICache.scala 96:32]
        tag1_16 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 56:28]
        tag1_16 <= tag1_31; // @[ICache.scala 56:28]
      end else begin
        tag1_16 <= _GEN_30;
      end
    end
    if (reset) begin // @[ICache.scala 49:26]
      tag1_17 <= 53'h0; // @[ICache.scala 49:26]
    end else if (5'h11 == index_addr) begin // @[ICache.scala 96:26]
      if (_block1_T) begin // @[ICache.scala 96:32]
        tag1_17 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 56:28]
        tag1_17 <= tag1_31; // @[ICache.scala 56:28]
      end else begin
        tag1_17 <= _GEN_30;
      end
    end
    if (reset) begin // @[ICache.scala 49:26]
      tag1_18 <= 53'h0; // @[ICache.scala 49:26]
    end else if (5'h12 == index_addr) begin // @[ICache.scala 96:26]
      if (_block1_T) begin // @[ICache.scala 96:32]
        tag1_18 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 56:28]
        tag1_18 <= tag1_31; // @[ICache.scala 56:28]
      end else begin
        tag1_18 <= _GEN_30;
      end
    end
    if (reset) begin // @[ICache.scala 49:26]
      tag1_19 <= 53'h0; // @[ICache.scala 49:26]
    end else if (5'h13 == index_addr) begin // @[ICache.scala 96:26]
      if (_block1_T) begin // @[ICache.scala 96:32]
        tag1_19 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 56:28]
        tag1_19 <= tag1_31; // @[ICache.scala 56:28]
      end else begin
        tag1_19 <= _GEN_30;
      end
    end
    if (reset) begin // @[ICache.scala 49:26]
      tag1_20 <= 53'h0; // @[ICache.scala 49:26]
    end else if (5'h14 == index_addr) begin // @[ICache.scala 96:26]
      if (_block1_T) begin // @[ICache.scala 96:32]
        tag1_20 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 56:28]
        tag1_20 <= tag1_31; // @[ICache.scala 56:28]
      end else begin
        tag1_20 <= _GEN_30;
      end
    end
    if (reset) begin // @[ICache.scala 49:26]
      tag1_21 <= 53'h0; // @[ICache.scala 49:26]
    end else if (5'h15 == index_addr) begin // @[ICache.scala 96:26]
      if (_block1_T) begin // @[ICache.scala 96:32]
        tag1_21 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 56:28]
        tag1_21 <= tag1_31; // @[ICache.scala 56:28]
      end else begin
        tag1_21 <= _GEN_30;
      end
    end
    if (reset) begin // @[ICache.scala 49:26]
      tag1_22 <= 53'h0; // @[ICache.scala 49:26]
    end else if (5'h16 == index_addr) begin // @[ICache.scala 96:26]
      if (_block1_T) begin // @[ICache.scala 96:32]
        tag1_22 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 56:28]
        tag1_22 <= tag1_31; // @[ICache.scala 56:28]
      end else begin
        tag1_22 <= _GEN_30;
      end
    end
    if (reset) begin // @[ICache.scala 49:26]
      tag1_23 <= 53'h0; // @[ICache.scala 49:26]
    end else if (5'h17 == index_addr) begin // @[ICache.scala 96:26]
      if (_block1_T) begin // @[ICache.scala 96:32]
        tag1_23 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 56:28]
        tag1_23 <= tag1_31; // @[ICache.scala 56:28]
      end else begin
        tag1_23 <= _GEN_30;
      end
    end
    if (reset) begin // @[ICache.scala 49:26]
      tag1_24 <= 53'h0; // @[ICache.scala 49:26]
    end else if (5'h18 == index_addr) begin // @[ICache.scala 96:26]
      if (_block1_T) begin // @[ICache.scala 96:32]
        tag1_24 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 56:28]
        tag1_24 <= tag1_31; // @[ICache.scala 56:28]
      end else begin
        tag1_24 <= _GEN_30;
      end
    end
    if (reset) begin // @[ICache.scala 49:26]
      tag1_25 <= 53'h0; // @[ICache.scala 49:26]
    end else if (5'h19 == index_addr) begin // @[ICache.scala 96:26]
      if (_block1_T) begin // @[ICache.scala 96:32]
        tag1_25 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 56:28]
        tag1_25 <= tag1_31; // @[ICache.scala 56:28]
      end else begin
        tag1_25 <= _GEN_30;
      end
    end
    if (reset) begin // @[ICache.scala 49:26]
      tag1_26 <= 53'h0; // @[ICache.scala 49:26]
    end else if (5'h1a == index_addr) begin // @[ICache.scala 96:26]
      if (_block1_T) begin // @[ICache.scala 96:32]
        tag1_26 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 56:28]
        tag1_26 <= tag1_31; // @[ICache.scala 56:28]
      end else begin
        tag1_26 <= _GEN_30;
      end
    end
    if (reset) begin // @[ICache.scala 49:26]
      tag1_27 <= 53'h0; // @[ICache.scala 49:26]
    end else if (5'h1b == index_addr) begin // @[ICache.scala 96:26]
      if (_block1_T) begin // @[ICache.scala 96:32]
        tag1_27 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 56:28]
        tag1_27 <= tag1_31; // @[ICache.scala 56:28]
      end else begin
        tag1_27 <= _GEN_30;
      end
    end
    if (reset) begin // @[ICache.scala 49:26]
      tag1_28 <= 53'h0; // @[ICache.scala 49:26]
    end else if (5'h1c == index_addr) begin // @[ICache.scala 96:26]
      if (_block1_T) begin // @[ICache.scala 96:32]
        tag1_28 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 56:28]
        tag1_28 <= tag1_31; // @[ICache.scala 56:28]
      end else begin
        tag1_28 <= _GEN_30;
      end
    end
    if (reset) begin // @[ICache.scala 49:26]
      tag1_29 <= 53'h0; // @[ICache.scala 49:26]
    end else if (5'h1d == index_addr) begin // @[ICache.scala 96:26]
      if (_block1_T) begin // @[ICache.scala 96:32]
        tag1_29 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 56:28]
        tag1_29 <= tag1_31; // @[ICache.scala 56:28]
      end else begin
        tag1_29 <= _GEN_30;
      end
    end
    if (reset) begin // @[ICache.scala 49:26]
      tag1_30 <= 53'h0; // @[ICache.scala 49:26]
    end else if (5'h1e == index_addr) begin // @[ICache.scala 96:26]
      if (_block1_T) begin // @[ICache.scala 96:32]
        tag1_30 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 56:28]
        tag1_30 <= tag1_31; // @[ICache.scala 56:28]
      end else begin
        tag1_30 <= _GEN_30;
      end
    end
    if (reset) begin // @[ICache.scala 49:26]
      tag1_31 <= 53'h0; // @[ICache.scala 49:26]
    end else if (5'h1f == index_addr) begin // @[ICache.scala 96:26]
      if (_block1_T) begin // @[ICache.scala 96:32]
        tag1_31 <= tag_addr;
      end else if (!(5'h1f == index_addr)) begin // @[ICache.scala 56:28]
        tag1_31 <= _GEN_30;
      end
    end
    if (reset) begin // @[ICache.scala 50:26]
      block1_0 <= 512'h0; // @[ICache.scala 50:26]
    end else if (5'h0 == index_addr) begin // @[ICache.scala 95:26]
      if (update & updateway1) begin // @[ICache.scala 95:32]
        block1_0 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 58:39]
        block1_0 <= block1_31; // @[ICache.scala 58:39]
      end else begin
        block1_0 <= _GEN_158;
      end
    end
    if (reset) begin // @[ICache.scala 50:26]
      block1_1 <= 512'h0; // @[ICache.scala 50:26]
    end else if (5'h1 == index_addr) begin // @[ICache.scala 95:26]
      if (update & updateway1) begin // @[ICache.scala 95:32]
        block1_1 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 58:39]
        block1_1 <= block1_31; // @[ICache.scala 58:39]
      end else begin
        block1_1 <= _GEN_158;
      end
    end
    if (reset) begin // @[ICache.scala 50:26]
      block1_2 <= 512'h0; // @[ICache.scala 50:26]
    end else if (5'h2 == index_addr) begin // @[ICache.scala 95:26]
      if (update & updateway1) begin // @[ICache.scala 95:32]
        block1_2 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 58:39]
        block1_2 <= block1_31; // @[ICache.scala 58:39]
      end else begin
        block1_2 <= _GEN_158;
      end
    end
    if (reset) begin // @[ICache.scala 50:26]
      block1_3 <= 512'h0; // @[ICache.scala 50:26]
    end else if (5'h3 == index_addr) begin // @[ICache.scala 95:26]
      if (update & updateway1) begin // @[ICache.scala 95:32]
        block1_3 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 58:39]
        block1_3 <= block1_31; // @[ICache.scala 58:39]
      end else begin
        block1_3 <= _GEN_158;
      end
    end
    if (reset) begin // @[ICache.scala 50:26]
      block1_4 <= 512'h0; // @[ICache.scala 50:26]
    end else if (5'h4 == index_addr) begin // @[ICache.scala 95:26]
      if (update & updateway1) begin // @[ICache.scala 95:32]
        block1_4 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 58:39]
        block1_4 <= block1_31; // @[ICache.scala 58:39]
      end else begin
        block1_4 <= _GEN_158;
      end
    end
    if (reset) begin // @[ICache.scala 50:26]
      block1_5 <= 512'h0; // @[ICache.scala 50:26]
    end else if (5'h5 == index_addr) begin // @[ICache.scala 95:26]
      if (update & updateway1) begin // @[ICache.scala 95:32]
        block1_5 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 58:39]
        block1_5 <= block1_31; // @[ICache.scala 58:39]
      end else begin
        block1_5 <= _GEN_158;
      end
    end
    if (reset) begin // @[ICache.scala 50:26]
      block1_6 <= 512'h0; // @[ICache.scala 50:26]
    end else if (5'h6 == index_addr) begin // @[ICache.scala 95:26]
      if (update & updateway1) begin // @[ICache.scala 95:32]
        block1_6 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 58:39]
        block1_6 <= block1_31; // @[ICache.scala 58:39]
      end else begin
        block1_6 <= _GEN_158;
      end
    end
    if (reset) begin // @[ICache.scala 50:26]
      block1_7 <= 512'h0; // @[ICache.scala 50:26]
    end else if (5'h7 == index_addr) begin // @[ICache.scala 95:26]
      if (update & updateway1) begin // @[ICache.scala 95:32]
        block1_7 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 58:39]
        block1_7 <= block1_31; // @[ICache.scala 58:39]
      end else begin
        block1_7 <= _GEN_158;
      end
    end
    if (reset) begin // @[ICache.scala 50:26]
      block1_8 <= 512'h0; // @[ICache.scala 50:26]
    end else if (5'h8 == index_addr) begin // @[ICache.scala 95:26]
      if (update & updateway1) begin // @[ICache.scala 95:32]
        block1_8 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 58:39]
        block1_8 <= block1_31; // @[ICache.scala 58:39]
      end else begin
        block1_8 <= _GEN_158;
      end
    end
    if (reset) begin // @[ICache.scala 50:26]
      block1_9 <= 512'h0; // @[ICache.scala 50:26]
    end else if (5'h9 == index_addr) begin // @[ICache.scala 95:26]
      if (update & updateway1) begin // @[ICache.scala 95:32]
        block1_9 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 58:39]
        block1_9 <= block1_31; // @[ICache.scala 58:39]
      end else begin
        block1_9 <= _GEN_158;
      end
    end
    if (reset) begin // @[ICache.scala 50:26]
      block1_10 <= 512'h0; // @[ICache.scala 50:26]
    end else if (5'ha == index_addr) begin // @[ICache.scala 95:26]
      if (update & updateway1) begin // @[ICache.scala 95:32]
        block1_10 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 58:39]
        block1_10 <= block1_31; // @[ICache.scala 58:39]
      end else begin
        block1_10 <= _GEN_158;
      end
    end
    if (reset) begin // @[ICache.scala 50:26]
      block1_11 <= 512'h0; // @[ICache.scala 50:26]
    end else if (5'hb == index_addr) begin // @[ICache.scala 95:26]
      if (update & updateway1) begin // @[ICache.scala 95:32]
        block1_11 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 58:39]
        block1_11 <= block1_31; // @[ICache.scala 58:39]
      end else begin
        block1_11 <= _GEN_158;
      end
    end
    if (reset) begin // @[ICache.scala 50:26]
      block1_12 <= 512'h0; // @[ICache.scala 50:26]
    end else if (5'hc == index_addr) begin // @[ICache.scala 95:26]
      if (update & updateway1) begin // @[ICache.scala 95:32]
        block1_12 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 58:39]
        block1_12 <= block1_31; // @[ICache.scala 58:39]
      end else begin
        block1_12 <= _GEN_158;
      end
    end
    if (reset) begin // @[ICache.scala 50:26]
      block1_13 <= 512'h0; // @[ICache.scala 50:26]
    end else if (5'hd == index_addr) begin // @[ICache.scala 95:26]
      if (update & updateway1) begin // @[ICache.scala 95:32]
        block1_13 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 58:39]
        block1_13 <= block1_31; // @[ICache.scala 58:39]
      end else begin
        block1_13 <= _GEN_158;
      end
    end
    if (reset) begin // @[ICache.scala 50:26]
      block1_14 <= 512'h0; // @[ICache.scala 50:26]
    end else if (5'he == index_addr) begin // @[ICache.scala 95:26]
      if (update & updateway1) begin // @[ICache.scala 95:32]
        block1_14 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 58:39]
        block1_14 <= block1_31; // @[ICache.scala 58:39]
      end else begin
        block1_14 <= _GEN_158;
      end
    end
    if (reset) begin // @[ICache.scala 50:26]
      block1_15 <= 512'h0; // @[ICache.scala 50:26]
    end else if (5'hf == index_addr) begin // @[ICache.scala 95:26]
      if (update & updateway1) begin // @[ICache.scala 95:32]
        block1_15 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 58:39]
        block1_15 <= block1_31; // @[ICache.scala 58:39]
      end else begin
        block1_15 <= _GEN_158;
      end
    end
    if (reset) begin // @[ICache.scala 50:26]
      block1_16 <= 512'h0; // @[ICache.scala 50:26]
    end else if (5'h10 == index_addr) begin // @[ICache.scala 95:26]
      if (update & updateway1) begin // @[ICache.scala 95:32]
        block1_16 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 58:39]
        block1_16 <= block1_31; // @[ICache.scala 58:39]
      end else begin
        block1_16 <= _GEN_158;
      end
    end
    if (reset) begin // @[ICache.scala 50:26]
      block1_17 <= 512'h0; // @[ICache.scala 50:26]
    end else if (5'h11 == index_addr) begin // @[ICache.scala 95:26]
      if (update & updateway1) begin // @[ICache.scala 95:32]
        block1_17 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 58:39]
        block1_17 <= block1_31; // @[ICache.scala 58:39]
      end else begin
        block1_17 <= _GEN_158;
      end
    end
    if (reset) begin // @[ICache.scala 50:26]
      block1_18 <= 512'h0; // @[ICache.scala 50:26]
    end else if (5'h12 == index_addr) begin // @[ICache.scala 95:26]
      if (update & updateway1) begin // @[ICache.scala 95:32]
        block1_18 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 58:39]
        block1_18 <= block1_31; // @[ICache.scala 58:39]
      end else begin
        block1_18 <= _GEN_158;
      end
    end
    if (reset) begin // @[ICache.scala 50:26]
      block1_19 <= 512'h0; // @[ICache.scala 50:26]
    end else if (5'h13 == index_addr) begin // @[ICache.scala 95:26]
      if (update & updateway1) begin // @[ICache.scala 95:32]
        block1_19 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 58:39]
        block1_19 <= block1_31; // @[ICache.scala 58:39]
      end else begin
        block1_19 <= _GEN_158;
      end
    end
    if (reset) begin // @[ICache.scala 50:26]
      block1_20 <= 512'h0; // @[ICache.scala 50:26]
    end else if (5'h14 == index_addr) begin // @[ICache.scala 95:26]
      if (update & updateway1) begin // @[ICache.scala 95:32]
        block1_20 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 58:39]
        block1_20 <= block1_31; // @[ICache.scala 58:39]
      end else begin
        block1_20 <= _GEN_158;
      end
    end
    if (reset) begin // @[ICache.scala 50:26]
      block1_21 <= 512'h0; // @[ICache.scala 50:26]
    end else if (5'h15 == index_addr) begin // @[ICache.scala 95:26]
      if (update & updateway1) begin // @[ICache.scala 95:32]
        block1_21 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 58:39]
        block1_21 <= block1_31; // @[ICache.scala 58:39]
      end else begin
        block1_21 <= _GEN_158;
      end
    end
    if (reset) begin // @[ICache.scala 50:26]
      block1_22 <= 512'h0; // @[ICache.scala 50:26]
    end else if (5'h16 == index_addr) begin // @[ICache.scala 95:26]
      if (update & updateway1) begin // @[ICache.scala 95:32]
        block1_22 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 58:39]
        block1_22 <= block1_31; // @[ICache.scala 58:39]
      end else begin
        block1_22 <= _GEN_158;
      end
    end
    if (reset) begin // @[ICache.scala 50:26]
      block1_23 <= 512'h0; // @[ICache.scala 50:26]
    end else if (5'h17 == index_addr) begin // @[ICache.scala 95:26]
      if (update & updateway1) begin // @[ICache.scala 95:32]
        block1_23 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 58:39]
        block1_23 <= block1_31; // @[ICache.scala 58:39]
      end else begin
        block1_23 <= _GEN_158;
      end
    end
    if (reset) begin // @[ICache.scala 50:26]
      block1_24 <= 512'h0; // @[ICache.scala 50:26]
    end else if (5'h18 == index_addr) begin // @[ICache.scala 95:26]
      if (update & updateway1) begin // @[ICache.scala 95:32]
        block1_24 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 58:39]
        block1_24 <= block1_31; // @[ICache.scala 58:39]
      end else begin
        block1_24 <= _GEN_158;
      end
    end
    if (reset) begin // @[ICache.scala 50:26]
      block1_25 <= 512'h0; // @[ICache.scala 50:26]
    end else if (5'h19 == index_addr) begin // @[ICache.scala 95:26]
      if (update & updateway1) begin // @[ICache.scala 95:32]
        block1_25 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 58:39]
        block1_25 <= block1_31; // @[ICache.scala 58:39]
      end else begin
        block1_25 <= _GEN_158;
      end
    end
    if (reset) begin // @[ICache.scala 50:26]
      block1_26 <= 512'h0; // @[ICache.scala 50:26]
    end else if (5'h1a == index_addr) begin // @[ICache.scala 95:26]
      if (update & updateway1) begin // @[ICache.scala 95:32]
        block1_26 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 58:39]
        block1_26 <= block1_31; // @[ICache.scala 58:39]
      end else begin
        block1_26 <= _GEN_158;
      end
    end
    if (reset) begin // @[ICache.scala 50:26]
      block1_27 <= 512'h0; // @[ICache.scala 50:26]
    end else if (5'h1b == index_addr) begin // @[ICache.scala 95:26]
      if (update & updateway1) begin // @[ICache.scala 95:32]
        block1_27 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 58:39]
        block1_27 <= block1_31; // @[ICache.scala 58:39]
      end else begin
        block1_27 <= _GEN_158;
      end
    end
    if (reset) begin // @[ICache.scala 50:26]
      block1_28 <= 512'h0; // @[ICache.scala 50:26]
    end else if (5'h1c == index_addr) begin // @[ICache.scala 95:26]
      if (update & updateway1) begin // @[ICache.scala 95:32]
        block1_28 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 58:39]
        block1_28 <= block1_31; // @[ICache.scala 58:39]
      end else begin
        block1_28 <= _GEN_158;
      end
    end
    if (reset) begin // @[ICache.scala 50:26]
      block1_29 <= 512'h0; // @[ICache.scala 50:26]
    end else if (5'h1d == index_addr) begin // @[ICache.scala 95:26]
      if (update & updateway1) begin // @[ICache.scala 95:32]
        block1_29 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 58:39]
        block1_29 <= block1_31; // @[ICache.scala 58:39]
      end else begin
        block1_29 <= _GEN_158;
      end
    end
    if (reset) begin // @[ICache.scala 50:26]
      block1_30 <= 512'h0; // @[ICache.scala 50:26]
    end else if (5'h1e == index_addr) begin // @[ICache.scala 95:26]
      if (update & updateway1) begin // @[ICache.scala 95:32]
        block1_30 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 58:39]
        block1_30 <= block1_31; // @[ICache.scala 58:39]
      end else begin
        block1_30 <= _GEN_158;
      end
    end
    if (reset) begin // @[ICache.scala 50:26]
      block1_31 <= 512'h0; // @[ICache.scala 50:26]
    end else if (5'h1f == index_addr) begin // @[ICache.scala 95:26]
      if (update & updateway1) begin // @[ICache.scala 95:32]
        block1_31 <= io_axi_data;
      end else if (!(5'h1f == index_addr)) begin // @[ICache.scala 58:39]
        block1_31 <= _GEN_158;
      end
    end
    if (reset) begin // @[ICache.scala 51:26]
      v2_0 <= 1'h0; // @[ICache.scala 51:26]
    end else if (5'h0 == index_addr) begin // @[ICache.scala 100:26]
      v2_0 <= _block2_T | _GEN_127; // @[ICache.scala 100:26]
    end
    if (reset) begin // @[ICache.scala 51:26]
      v2_1 <= 1'h0; // @[ICache.scala 51:26]
    end else if (5'h1 == index_addr) begin // @[ICache.scala 100:26]
      v2_1 <= _block2_T | _GEN_127; // @[ICache.scala 100:26]
    end
    if (reset) begin // @[ICache.scala 51:26]
      v2_2 <= 1'h0; // @[ICache.scala 51:26]
    end else if (5'h2 == index_addr) begin // @[ICache.scala 100:26]
      v2_2 <= _block2_T | _GEN_127; // @[ICache.scala 100:26]
    end
    if (reset) begin // @[ICache.scala 51:26]
      v2_3 <= 1'h0; // @[ICache.scala 51:26]
    end else if (5'h3 == index_addr) begin // @[ICache.scala 100:26]
      v2_3 <= _block2_T | _GEN_127; // @[ICache.scala 100:26]
    end
    if (reset) begin // @[ICache.scala 51:26]
      v2_4 <= 1'h0; // @[ICache.scala 51:26]
    end else if (5'h4 == index_addr) begin // @[ICache.scala 100:26]
      v2_4 <= _block2_T | _GEN_127; // @[ICache.scala 100:26]
    end
    if (reset) begin // @[ICache.scala 51:26]
      v2_5 <= 1'h0; // @[ICache.scala 51:26]
    end else if (5'h5 == index_addr) begin // @[ICache.scala 100:26]
      v2_5 <= _block2_T | _GEN_127; // @[ICache.scala 100:26]
    end
    if (reset) begin // @[ICache.scala 51:26]
      v2_6 <= 1'h0; // @[ICache.scala 51:26]
    end else if (5'h6 == index_addr) begin // @[ICache.scala 100:26]
      v2_6 <= _block2_T | _GEN_127; // @[ICache.scala 100:26]
    end
    if (reset) begin // @[ICache.scala 51:26]
      v2_7 <= 1'h0; // @[ICache.scala 51:26]
    end else if (5'h7 == index_addr) begin // @[ICache.scala 100:26]
      v2_7 <= _block2_T | _GEN_127; // @[ICache.scala 100:26]
    end
    if (reset) begin // @[ICache.scala 51:26]
      v2_8 <= 1'h0; // @[ICache.scala 51:26]
    end else if (5'h8 == index_addr) begin // @[ICache.scala 100:26]
      v2_8 <= _block2_T | _GEN_127; // @[ICache.scala 100:26]
    end
    if (reset) begin // @[ICache.scala 51:26]
      v2_9 <= 1'h0; // @[ICache.scala 51:26]
    end else if (5'h9 == index_addr) begin // @[ICache.scala 100:26]
      v2_9 <= _block2_T | _GEN_127; // @[ICache.scala 100:26]
    end
    if (reset) begin // @[ICache.scala 51:26]
      v2_10 <= 1'h0; // @[ICache.scala 51:26]
    end else if (5'ha == index_addr) begin // @[ICache.scala 100:26]
      v2_10 <= _block2_T | _GEN_127; // @[ICache.scala 100:26]
    end
    if (reset) begin // @[ICache.scala 51:26]
      v2_11 <= 1'h0; // @[ICache.scala 51:26]
    end else if (5'hb == index_addr) begin // @[ICache.scala 100:26]
      v2_11 <= _block2_T | _GEN_127; // @[ICache.scala 100:26]
    end
    if (reset) begin // @[ICache.scala 51:26]
      v2_12 <= 1'h0; // @[ICache.scala 51:26]
    end else if (5'hc == index_addr) begin // @[ICache.scala 100:26]
      v2_12 <= _block2_T | _GEN_127; // @[ICache.scala 100:26]
    end
    if (reset) begin // @[ICache.scala 51:26]
      v2_13 <= 1'h0; // @[ICache.scala 51:26]
    end else if (5'hd == index_addr) begin // @[ICache.scala 100:26]
      v2_13 <= _block2_T | _GEN_127; // @[ICache.scala 100:26]
    end
    if (reset) begin // @[ICache.scala 51:26]
      v2_14 <= 1'h0; // @[ICache.scala 51:26]
    end else if (5'he == index_addr) begin // @[ICache.scala 100:26]
      v2_14 <= _block2_T | _GEN_127; // @[ICache.scala 100:26]
    end
    if (reset) begin // @[ICache.scala 51:26]
      v2_15 <= 1'h0; // @[ICache.scala 51:26]
    end else if (5'hf == index_addr) begin // @[ICache.scala 100:26]
      v2_15 <= _block2_T | _GEN_127; // @[ICache.scala 100:26]
    end
    if (reset) begin // @[ICache.scala 51:26]
      v2_16 <= 1'h0; // @[ICache.scala 51:26]
    end else if (5'h10 == index_addr) begin // @[ICache.scala 100:26]
      v2_16 <= _block2_T | _GEN_127; // @[ICache.scala 100:26]
    end
    if (reset) begin // @[ICache.scala 51:26]
      v2_17 <= 1'h0; // @[ICache.scala 51:26]
    end else if (5'h11 == index_addr) begin // @[ICache.scala 100:26]
      v2_17 <= _block2_T | _GEN_127; // @[ICache.scala 100:26]
    end
    if (reset) begin // @[ICache.scala 51:26]
      v2_18 <= 1'h0; // @[ICache.scala 51:26]
    end else if (5'h12 == index_addr) begin // @[ICache.scala 100:26]
      v2_18 <= _block2_T | _GEN_127; // @[ICache.scala 100:26]
    end
    if (reset) begin // @[ICache.scala 51:26]
      v2_19 <= 1'h0; // @[ICache.scala 51:26]
    end else if (5'h13 == index_addr) begin // @[ICache.scala 100:26]
      v2_19 <= _block2_T | _GEN_127; // @[ICache.scala 100:26]
    end
    if (reset) begin // @[ICache.scala 51:26]
      v2_20 <= 1'h0; // @[ICache.scala 51:26]
    end else if (5'h14 == index_addr) begin // @[ICache.scala 100:26]
      v2_20 <= _block2_T | _GEN_127; // @[ICache.scala 100:26]
    end
    if (reset) begin // @[ICache.scala 51:26]
      v2_21 <= 1'h0; // @[ICache.scala 51:26]
    end else if (5'h15 == index_addr) begin // @[ICache.scala 100:26]
      v2_21 <= _block2_T | _GEN_127; // @[ICache.scala 100:26]
    end
    if (reset) begin // @[ICache.scala 51:26]
      v2_22 <= 1'h0; // @[ICache.scala 51:26]
    end else if (5'h16 == index_addr) begin // @[ICache.scala 100:26]
      v2_22 <= _block2_T | _GEN_127; // @[ICache.scala 100:26]
    end
    if (reset) begin // @[ICache.scala 51:26]
      v2_23 <= 1'h0; // @[ICache.scala 51:26]
    end else if (5'h17 == index_addr) begin // @[ICache.scala 100:26]
      v2_23 <= _block2_T | _GEN_127; // @[ICache.scala 100:26]
    end
    if (reset) begin // @[ICache.scala 51:26]
      v2_24 <= 1'h0; // @[ICache.scala 51:26]
    end else if (5'h18 == index_addr) begin // @[ICache.scala 100:26]
      v2_24 <= _block2_T | _GEN_127; // @[ICache.scala 100:26]
    end
    if (reset) begin // @[ICache.scala 51:26]
      v2_25 <= 1'h0; // @[ICache.scala 51:26]
    end else if (5'h19 == index_addr) begin // @[ICache.scala 100:26]
      v2_25 <= _block2_T | _GEN_127; // @[ICache.scala 100:26]
    end
    if (reset) begin // @[ICache.scala 51:26]
      v2_26 <= 1'h0; // @[ICache.scala 51:26]
    end else if (5'h1a == index_addr) begin // @[ICache.scala 100:26]
      v2_26 <= _block2_T | _GEN_127; // @[ICache.scala 100:26]
    end
    if (reset) begin // @[ICache.scala 51:26]
      v2_27 <= 1'h0; // @[ICache.scala 51:26]
    end else if (5'h1b == index_addr) begin // @[ICache.scala 100:26]
      v2_27 <= _block2_T | _GEN_127; // @[ICache.scala 100:26]
    end
    if (reset) begin // @[ICache.scala 51:26]
      v2_28 <= 1'h0; // @[ICache.scala 51:26]
    end else if (5'h1c == index_addr) begin // @[ICache.scala 100:26]
      v2_28 <= _block2_T | _GEN_127; // @[ICache.scala 100:26]
    end
    if (reset) begin // @[ICache.scala 51:26]
      v2_29 <= 1'h0; // @[ICache.scala 51:26]
    end else if (5'h1d == index_addr) begin // @[ICache.scala 100:26]
      v2_29 <= _block2_T | _GEN_127; // @[ICache.scala 100:26]
    end
    if (reset) begin // @[ICache.scala 51:26]
      v2_30 <= 1'h0; // @[ICache.scala 51:26]
    end else if (5'h1e == index_addr) begin // @[ICache.scala 100:26]
      v2_30 <= _block2_T | _GEN_127; // @[ICache.scala 100:26]
    end
    if (reset) begin // @[ICache.scala 51:26]
      v2_31 <= 1'h0; // @[ICache.scala 51:26]
    end else if (5'h1f == index_addr) begin // @[ICache.scala 100:26]
      v2_31 <= _block2_T | _GEN_127; // @[ICache.scala 100:26]
    end
    if (reset) begin // @[ICache.scala 52:26]
      age2_0 <= 1'h0; // @[ICache.scala 52:26]
    end else if (5'h0 == index_addr) begin // @[ICache.scala 67:22]
      if (_age1_T) begin // @[ICache.scala 67:28]
        age2_0 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 67:28]
        age2_0 <= age2_31; // @[ICache.scala 67:28]
      end else begin
        age2_0 <= _GEN_286;
      end
    end
    if (reset) begin // @[ICache.scala 52:26]
      age2_1 <= 1'h0; // @[ICache.scala 52:26]
    end else if (5'h1 == index_addr) begin // @[ICache.scala 67:22]
      if (_age1_T) begin // @[ICache.scala 67:28]
        age2_1 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 67:28]
        age2_1 <= age2_31; // @[ICache.scala 67:28]
      end else begin
        age2_1 <= _GEN_286;
      end
    end
    if (reset) begin // @[ICache.scala 52:26]
      age2_2 <= 1'h0; // @[ICache.scala 52:26]
    end else if (5'h2 == index_addr) begin // @[ICache.scala 67:22]
      if (_age1_T) begin // @[ICache.scala 67:28]
        age2_2 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 67:28]
        age2_2 <= age2_31; // @[ICache.scala 67:28]
      end else begin
        age2_2 <= _GEN_286;
      end
    end
    if (reset) begin // @[ICache.scala 52:26]
      age2_3 <= 1'h0; // @[ICache.scala 52:26]
    end else if (5'h3 == index_addr) begin // @[ICache.scala 67:22]
      if (_age1_T) begin // @[ICache.scala 67:28]
        age2_3 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 67:28]
        age2_3 <= age2_31; // @[ICache.scala 67:28]
      end else begin
        age2_3 <= _GEN_286;
      end
    end
    if (reset) begin // @[ICache.scala 52:26]
      age2_4 <= 1'h0; // @[ICache.scala 52:26]
    end else if (5'h4 == index_addr) begin // @[ICache.scala 67:22]
      if (_age1_T) begin // @[ICache.scala 67:28]
        age2_4 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 67:28]
        age2_4 <= age2_31; // @[ICache.scala 67:28]
      end else begin
        age2_4 <= _GEN_286;
      end
    end
    if (reset) begin // @[ICache.scala 52:26]
      age2_5 <= 1'h0; // @[ICache.scala 52:26]
    end else if (5'h5 == index_addr) begin // @[ICache.scala 67:22]
      if (_age1_T) begin // @[ICache.scala 67:28]
        age2_5 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 67:28]
        age2_5 <= age2_31; // @[ICache.scala 67:28]
      end else begin
        age2_5 <= _GEN_286;
      end
    end
    if (reset) begin // @[ICache.scala 52:26]
      age2_6 <= 1'h0; // @[ICache.scala 52:26]
    end else if (5'h6 == index_addr) begin // @[ICache.scala 67:22]
      if (_age1_T) begin // @[ICache.scala 67:28]
        age2_6 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 67:28]
        age2_6 <= age2_31; // @[ICache.scala 67:28]
      end else begin
        age2_6 <= _GEN_286;
      end
    end
    if (reset) begin // @[ICache.scala 52:26]
      age2_7 <= 1'h0; // @[ICache.scala 52:26]
    end else if (5'h7 == index_addr) begin // @[ICache.scala 67:22]
      if (_age1_T) begin // @[ICache.scala 67:28]
        age2_7 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 67:28]
        age2_7 <= age2_31; // @[ICache.scala 67:28]
      end else begin
        age2_7 <= _GEN_286;
      end
    end
    if (reset) begin // @[ICache.scala 52:26]
      age2_8 <= 1'h0; // @[ICache.scala 52:26]
    end else if (5'h8 == index_addr) begin // @[ICache.scala 67:22]
      if (_age1_T) begin // @[ICache.scala 67:28]
        age2_8 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 67:28]
        age2_8 <= age2_31; // @[ICache.scala 67:28]
      end else begin
        age2_8 <= _GEN_286;
      end
    end
    if (reset) begin // @[ICache.scala 52:26]
      age2_9 <= 1'h0; // @[ICache.scala 52:26]
    end else if (5'h9 == index_addr) begin // @[ICache.scala 67:22]
      if (_age1_T) begin // @[ICache.scala 67:28]
        age2_9 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 67:28]
        age2_9 <= age2_31; // @[ICache.scala 67:28]
      end else begin
        age2_9 <= _GEN_286;
      end
    end
    if (reset) begin // @[ICache.scala 52:26]
      age2_10 <= 1'h0; // @[ICache.scala 52:26]
    end else if (5'ha == index_addr) begin // @[ICache.scala 67:22]
      if (_age1_T) begin // @[ICache.scala 67:28]
        age2_10 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 67:28]
        age2_10 <= age2_31; // @[ICache.scala 67:28]
      end else begin
        age2_10 <= _GEN_286;
      end
    end
    if (reset) begin // @[ICache.scala 52:26]
      age2_11 <= 1'h0; // @[ICache.scala 52:26]
    end else if (5'hb == index_addr) begin // @[ICache.scala 67:22]
      if (_age1_T) begin // @[ICache.scala 67:28]
        age2_11 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 67:28]
        age2_11 <= age2_31; // @[ICache.scala 67:28]
      end else begin
        age2_11 <= _GEN_286;
      end
    end
    if (reset) begin // @[ICache.scala 52:26]
      age2_12 <= 1'h0; // @[ICache.scala 52:26]
    end else if (5'hc == index_addr) begin // @[ICache.scala 67:22]
      if (_age1_T) begin // @[ICache.scala 67:28]
        age2_12 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 67:28]
        age2_12 <= age2_31; // @[ICache.scala 67:28]
      end else begin
        age2_12 <= _GEN_286;
      end
    end
    if (reset) begin // @[ICache.scala 52:26]
      age2_13 <= 1'h0; // @[ICache.scala 52:26]
    end else if (5'hd == index_addr) begin // @[ICache.scala 67:22]
      if (_age1_T) begin // @[ICache.scala 67:28]
        age2_13 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 67:28]
        age2_13 <= age2_31; // @[ICache.scala 67:28]
      end else begin
        age2_13 <= _GEN_286;
      end
    end
    if (reset) begin // @[ICache.scala 52:26]
      age2_14 <= 1'h0; // @[ICache.scala 52:26]
    end else if (5'he == index_addr) begin // @[ICache.scala 67:22]
      if (_age1_T) begin // @[ICache.scala 67:28]
        age2_14 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 67:28]
        age2_14 <= age2_31; // @[ICache.scala 67:28]
      end else begin
        age2_14 <= _GEN_286;
      end
    end
    if (reset) begin // @[ICache.scala 52:26]
      age2_15 <= 1'h0; // @[ICache.scala 52:26]
    end else if (5'hf == index_addr) begin // @[ICache.scala 67:22]
      if (_age1_T) begin // @[ICache.scala 67:28]
        age2_15 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 67:28]
        age2_15 <= age2_31; // @[ICache.scala 67:28]
      end else begin
        age2_15 <= _GEN_286;
      end
    end
    if (reset) begin // @[ICache.scala 52:26]
      age2_16 <= 1'h0; // @[ICache.scala 52:26]
    end else if (5'h10 == index_addr) begin // @[ICache.scala 67:22]
      if (_age1_T) begin // @[ICache.scala 67:28]
        age2_16 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 67:28]
        age2_16 <= age2_31; // @[ICache.scala 67:28]
      end else begin
        age2_16 <= _GEN_286;
      end
    end
    if (reset) begin // @[ICache.scala 52:26]
      age2_17 <= 1'h0; // @[ICache.scala 52:26]
    end else if (5'h11 == index_addr) begin // @[ICache.scala 67:22]
      if (_age1_T) begin // @[ICache.scala 67:28]
        age2_17 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 67:28]
        age2_17 <= age2_31; // @[ICache.scala 67:28]
      end else begin
        age2_17 <= _GEN_286;
      end
    end
    if (reset) begin // @[ICache.scala 52:26]
      age2_18 <= 1'h0; // @[ICache.scala 52:26]
    end else if (5'h12 == index_addr) begin // @[ICache.scala 67:22]
      if (_age1_T) begin // @[ICache.scala 67:28]
        age2_18 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 67:28]
        age2_18 <= age2_31; // @[ICache.scala 67:28]
      end else begin
        age2_18 <= _GEN_286;
      end
    end
    if (reset) begin // @[ICache.scala 52:26]
      age2_19 <= 1'h0; // @[ICache.scala 52:26]
    end else if (5'h13 == index_addr) begin // @[ICache.scala 67:22]
      if (_age1_T) begin // @[ICache.scala 67:28]
        age2_19 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 67:28]
        age2_19 <= age2_31; // @[ICache.scala 67:28]
      end else begin
        age2_19 <= _GEN_286;
      end
    end
    if (reset) begin // @[ICache.scala 52:26]
      age2_20 <= 1'h0; // @[ICache.scala 52:26]
    end else if (5'h14 == index_addr) begin // @[ICache.scala 67:22]
      if (_age1_T) begin // @[ICache.scala 67:28]
        age2_20 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 67:28]
        age2_20 <= age2_31; // @[ICache.scala 67:28]
      end else begin
        age2_20 <= _GEN_286;
      end
    end
    if (reset) begin // @[ICache.scala 52:26]
      age2_21 <= 1'h0; // @[ICache.scala 52:26]
    end else if (5'h15 == index_addr) begin // @[ICache.scala 67:22]
      if (_age1_T) begin // @[ICache.scala 67:28]
        age2_21 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 67:28]
        age2_21 <= age2_31; // @[ICache.scala 67:28]
      end else begin
        age2_21 <= _GEN_286;
      end
    end
    if (reset) begin // @[ICache.scala 52:26]
      age2_22 <= 1'h0; // @[ICache.scala 52:26]
    end else if (5'h16 == index_addr) begin // @[ICache.scala 67:22]
      if (_age1_T) begin // @[ICache.scala 67:28]
        age2_22 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 67:28]
        age2_22 <= age2_31; // @[ICache.scala 67:28]
      end else begin
        age2_22 <= _GEN_286;
      end
    end
    if (reset) begin // @[ICache.scala 52:26]
      age2_23 <= 1'h0; // @[ICache.scala 52:26]
    end else if (5'h17 == index_addr) begin // @[ICache.scala 67:22]
      if (_age1_T) begin // @[ICache.scala 67:28]
        age2_23 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 67:28]
        age2_23 <= age2_31; // @[ICache.scala 67:28]
      end else begin
        age2_23 <= _GEN_286;
      end
    end
    if (reset) begin // @[ICache.scala 52:26]
      age2_24 <= 1'h0; // @[ICache.scala 52:26]
    end else if (5'h18 == index_addr) begin // @[ICache.scala 67:22]
      if (_age1_T) begin // @[ICache.scala 67:28]
        age2_24 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 67:28]
        age2_24 <= age2_31; // @[ICache.scala 67:28]
      end else begin
        age2_24 <= _GEN_286;
      end
    end
    if (reset) begin // @[ICache.scala 52:26]
      age2_25 <= 1'h0; // @[ICache.scala 52:26]
    end else if (5'h19 == index_addr) begin // @[ICache.scala 67:22]
      if (_age1_T) begin // @[ICache.scala 67:28]
        age2_25 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 67:28]
        age2_25 <= age2_31; // @[ICache.scala 67:28]
      end else begin
        age2_25 <= _GEN_286;
      end
    end
    if (reset) begin // @[ICache.scala 52:26]
      age2_26 <= 1'h0; // @[ICache.scala 52:26]
    end else if (5'h1a == index_addr) begin // @[ICache.scala 67:22]
      if (_age1_T) begin // @[ICache.scala 67:28]
        age2_26 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 67:28]
        age2_26 <= age2_31; // @[ICache.scala 67:28]
      end else begin
        age2_26 <= _GEN_286;
      end
    end
    if (reset) begin // @[ICache.scala 52:26]
      age2_27 <= 1'h0; // @[ICache.scala 52:26]
    end else if (5'h1b == index_addr) begin // @[ICache.scala 67:22]
      if (_age1_T) begin // @[ICache.scala 67:28]
        age2_27 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 67:28]
        age2_27 <= age2_31; // @[ICache.scala 67:28]
      end else begin
        age2_27 <= _GEN_286;
      end
    end
    if (reset) begin // @[ICache.scala 52:26]
      age2_28 <= 1'h0; // @[ICache.scala 52:26]
    end else if (5'h1c == index_addr) begin // @[ICache.scala 67:22]
      if (_age1_T) begin // @[ICache.scala 67:28]
        age2_28 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 67:28]
        age2_28 <= age2_31; // @[ICache.scala 67:28]
      end else begin
        age2_28 <= _GEN_286;
      end
    end
    if (reset) begin // @[ICache.scala 52:26]
      age2_29 <= 1'h0; // @[ICache.scala 52:26]
    end else if (5'h1d == index_addr) begin // @[ICache.scala 67:22]
      if (_age1_T) begin // @[ICache.scala 67:28]
        age2_29 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 67:28]
        age2_29 <= age2_31; // @[ICache.scala 67:28]
      end else begin
        age2_29 <= _GEN_286;
      end
    end
    if (reset) begin // @[ICache.scala 52:26]
      age2_30 <= 1'h0; // @[ICache.scala 52:26]
    end else if (5'h1e == index_addr) begin // @[ICache.scala 67:22]
      if (_age1_T) begin // @[ICache.scala 67:28]
        age2_30 <= hit2;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 67:28]
        age2_30 <= age2_31; // @[ICache.scala 67:28]
      end else begin
        age2_30 <= _GEN_286;
      end
    end
    if (reset) begin // @[ICache.scala 52:26]
      age2_31 <= 1'h0; // @[ICache.scala 52:26]
    end else if (5'h1f == index_addr) begin // @[ICache.scala 67:22]
      if (_age1_T) begin // @[ICache.scala 67:28]
        age2_31 <= hit2;
      end else if (!(5'h1f == index_addr)) begin // @[ICache.scala 67:28]
        age2_31 <= _GEN_286;
      end
    end
    if (reset) begin // @[ICache.scala 53:26]
      tag2_0 <= 53'h0; // @[ICache.scala 53:26]
    end else if (5'h0 == index_addr) begin // @[ICache.scala 99:26]
      if (_block2_T) begin // @[ICache.scala 99:32]
        tag2_0 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 57:28]
        tag2_0 <= tag2_31; // @[ICache.scala 57:28]
      end else begin
        tag2_0 <= _GEN_94;
      end
    end
    if (reset) begin // @[ICache.scala 53:26]
      tag2_1 <= 53'h0; // @[ICache.scala 53:26]
    end else if (5'h1 == index_addr) begin // @[ICache.scala 99:26]
      if (_block2_T) begin // @[ICache.scala 99:32]
        tag2_1 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 57:28]
        tag2_1 <= tag2_31; // @[ICache.scala 57:28]
      end else begin
        tag2_1 <= _GEN_94;
      end
    end
    if (reset) begin // @[ICache.scala 53:26]
      tag2_2 <= 53'h0; // @[ICache.scala 53:26]
    end else if (5'h2 == index_addr) begin // @[ICache.scala 99:26]
      if (_block2_T) begin // @[ICache.scala 99:32]
        tag2_2 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 57:28]
        tag2_2 <= tag2_31; // @[ICache.scala 57:28]
      end else begin
        tag2_2 <= _GEN_94;
      end
    end
    if (reset) begin // @[ICache.scala 53:26]
      tag2_3 <= 53'h0; // @[ICache.scala 53:26]
    end else if (5'h3 == index_addr) begin // @[ICache.scala 99:26]
      if (_block2_T) begin // @[ICache.scala 99:32]
        tag2_3 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 57:28]
        tag2_3 <= tag2_31; // @[ICache.scala 57:28]
      end else begin
        tag2_3 <= _GEN_94;
      end
    end
    if (reset) begin // @[ICache.scala 53:26]
      tag2_4 <= 53'h0; // @[ICache.scala 53:26]
    end else if (5'h4 == index_addr) begin // @[ICache.scala 99:26]
      if (_block2_T) begin // @[ICache.scala 99:32]
        tag2_4 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 57:28]
        tag2_4 <= tag2_31; // @[ICache.scala 57:28]
      end else begin
        tag2_4 <= _GEN_94;
      end
    end
    if (reset) begin // @[ICache.scala 53:26]
      tag2_5 <= 53'h0; // @[ICache.scala 53:26]
    end else if (5'h5 == index_addr) begin // @[ICache.scala 99:26]
      if (_block2_T) begin // @[ICache.scala 99:32]
        tag2_5 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 57:28]
        tag2_5 <= tag2_31; // @[ICache.scala 57:28]
      end else begin
        tag2_5 <= _GEN_94;
      end
    end
    if (reset) begin // @[ICache.scala 53:26]
      tag2_6 <= 53'h0; // @[ICache.scala 53:26]
    end else if (5'h6 == index_addr) begin // @[ICache.scala 99:26]
      if (_block2_T) begin // @[ICache.scala 99:32]
        tag2_6 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 57:28]
        tag2_6 <= tag2_31; // @[ICache.scala 57:28]
      end else begin
        tag2_6 <= _GEN_94;
      end
    end
    if (reset) begin // @[ICache.scala 53:26]
      tag2_7 <= 53'h0; // @[ICache.scala 53:26]
    end else if (5'h7 == index_addr) begin // @[ICache.scala 99:26]
      if (_block2_T) begin // @[ICache.scala 99:32]
        tag2_7 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 57:28]
        tag2_7 <= tag2_31; // @[ICache.scala 57:28]
      end else begin
        tag2_7 <= _GEN_94;
      end
    end
    if (reset) begin // @[ICache.scala 53:26]
      tag2_8 <= 53'h0; // @[ICache.scala 53:26]
    end else if (5'h8 == index_addr) begin // @[ICache.scala 99:26]
      if (_block2_T) begin // @[ICache.scala 99:32]
        tag2_8 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 57:28]
        tag2_8 <= tag2_31; // @[ICache.scala 57:28]
      end else begin
        tag2_8 <= _GEN_94;
      end
    end
    if (reset) begin // @[ICache.scala 53:26]
      tag2_9 <= 53'h0; // @[ICache.scala 53:26]
    end else if (5'h9 == index_addr) begin // @[ICache.scala 99:26]
      if (_block2_T) begin // @[ICache.scala 99:32]
        tag2_9 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 57:28]
        tag2_9 <= tag2_31; // @[ICache.scala 57:28]
      end else begin
        tag2_9 <= _GEN_94;
      end
    end
    if (reset) begin // @[ICache.scala 53:26]
      tag2_10 <= 53'h0; // @[ICache.scala 53:26]
    end else if (5'ha == index_addr) begin // @[ICache.scala 99:26]
      if (_block2_T) begin // @[ICache.scala 99:32]
        tag2_10 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 57:28]
        tag2_10 <= tag2_31; // @[ICache.scala 57:28]
      end else begin
        tag2_10 <= _GEN_94;
      end
    end
    if (reset) begin // @[ICache.scala 53:26]
      tag2_11 <= 53'h0; // @[ICache.scala 53:26]
    end else if (5'hb == index_addr) begin // @[ICache.scala 99:26]
      if (_block2_T) begin // @[ICache.scala 99:32]
        tag2_11 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 57:28]
        tag2_11 <= tag2_31; // @[ICache.scala 57:28]
      end else begin
        tag2_11 <= _GEN_94;
      end
    end
    if (reset) begin // @[ICache.scala 53:26]
      tag2_12 <= 53'h0; // @[ICache.scala 53:26]
    end else if (5'hc == index_addr) begin // @[ICache.scala 99:26]
      if (_block2_T) begin // @[ICache.scala 99:32]
        tag2_12 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 57:28]
        tag2_12 <= tag2_31; // @[ICache.scala 57:28]
      end else begin
        tag2_12 <= _GEN_94;
      end
    end
    if (reset) begin // @[ICache.scala 53:26]
      tag2_13 <= 53'h0; // @[ICache.scala 53:26]
    end else if (5'hd == index_addr) begin // @[ICache.scala 99:26]
      if (_block2_T) begin // @[ICache.scala 99:32]
        tag2_13 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 57:28]
        tag2_13 <= tag2_31; // @[ICache.scala 57:28]
      end else begin
        tag2_13 <= _GEN_94;
      end
    end
    if (reset) begin // @[ICache.scala 53:26]
      tag2_14 <= 53'h0; // @[ICache.scala 53:26]
    end else if (5'he == index_addr) begin // @[ICache.scala 99:26]
      if (_block2_T) begin // @[ICache.scala 99:32]
        tag2_14 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 57:28]
        tag2_14 <= tag2_31; // @[ICache.scala 57:28]
      end else begin
        tag2_14 <= _GEN_94;
      end
    end
    if (reset) begin // @[ICache.scala 53:26]
      tag2_15 <= 53'h0; // @[ICache.scala 53:26]
    end else if (5'hf == index_addr) begin // @[ICache.scala 99:26]
      if (_block2_T) begin // @[ICache.scala 99:32]
        tag2_15 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 57:28]
        tag2_15 <= tag2_31; // @[ICache.scala 57:28]
      end else begin
        tag2_15 <= _GEN_94;
      end
    end
    if (reset) begin // @[ICache.scala 53:26]
      tag2_16 <= 53'h0; // @[ICache.scala 53:26]
    end else if (5'h10 == index_addr) begin // @[ICache.scala 99:26]
      if (_block2_T) begin // @[ICache.scala 99:32]
        tag2_16 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 57:28]
        tag2_16 <= tag2_31; // @[ICache.scala 57:28]
      end else begin
        tag2_16 <= _GEN_94;
      end
    end
    if (reset) begin // @[ICache.scala 53:26]
      tag2_17 <= 53'h0; // @[ICache.scala 53:26]
    end else if (5'h11 == index_addr) begin // @[ICache.scala 99:26]
      if (_block2_T) begin // @[ICache.scala 99:32]
        tag2_17 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 57:28]
        tag2_17 <= tag2_31; // @[ICache.scala 57:28]
      end else begin
        tag2_17 <= _GEN_94;
      end
    end
    if (reset) begin // @[ICache.scala 53:26]
      tag2_18 <= 53'h0; // @[ICache.scala 53:26]
    end else if (5'h12 == index_addr) begin // @[ICache.scala 99:26]
      if (_block2_T) begin // @[ICache.scala 99:32]
        tag2_18 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 57:28]
        tag2_18 <= tag2_31; // @[ICache.scala 57:28]
      end else begin
        tag2_18 <= _GEN_94;
      end
    end
    if (reset) begin // @[ICache.scala 53:26]
      tag2_19 <= 53'h0; // @[ICache.scala 53:26]
    end else if (5'h13 == index_addr) begin // @[ICache.scala 99:26]
      if (_block2_T) begin // @[ICache.scala 99:32]
        tag2_19 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 57:28]
        tag2_19 <= tag2_31; // @[ICache.scala 57:28]
      end else begin
        tag2_19 <= _GEN_94;
      end
    end
    if (reset) begin // @[ICache.scala 53:26]
      tag2_20 <= 53'h0; // @[ICache.scala 53:26]
    end else if (5'h14 == index_addr) begin // @[ICache.scala 99:26]
      if (_block2_T) begin // @[ICache.scala 99:32]
        tag2_20 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 57:28]
        tag2_20 <= tag2_31; // @[ICache.scala 57:28]
      end else begin
        tag2_20 <= _GEN_94;
      end
    end
    if (reset) begin // @[ICache.scala 53:26]
      tag2_21 <= 53'h0; // @[ICache.scala 53:26]
    end else if (5'h15 == index_addr) begin // @[ICache.scala 99:26]
      if (_block2_T) begin // @[ICache.scala 99:32]
        tag2_21 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 57:28]
        tag2_21 <= tag2_31; // @[ICache.scala 57:28]
      end else begin
        tag2_21 <= _GEN_94;
      end
    end
    if (reset) begin // @[ICache.scala 53:26]
      tag2_22 <= 53'h0; // @[ICache.scala 53:26]
    end else if (5'h16 == index_addr) begin // @[ICache.scala 99:26]
      if (_block2_T) begin // @[ICache.scala 99:32]
        tag2_22 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 57:28]
        tag2_22 <= tag2_31; // @[ICache.scala 57:28]
      end else begin
        tag2_22 <= _GEN_94;
      end
    end
    if (reset) begin // @[ICache.scala 53:26]
      tag2_23 <= 53'h0; // @[ICache.scala 53:26]
    end else if (5'h17 == index_addr) begin // @[ICache.scala 99:26]
      if (_block2_T) begin // @[ICache.scala 99:32]
        tag2_23 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 57:28]
        tag2_23 <= tag2_31; // @[ICache.scala 57:28]
      end else begin
        tag2_23 <= _GEN_94;
      end
    end
    if (reset) begin // @[ICache.scala 53:26]
      tag2_24 <= 53'h0; // @[ICache.scala 53:26]
    end else if (5'h18 == index_addr) begin // @[ICache.scala 99:26]
      if (_block2_T) begin // @[ICache.scala 99:32]
        tag2_24 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 57:28]
        tag2_24 <= tag2_31; // @[ICache.scala 57:28]
      end else begin
        tag2_24 <= _GEN_94;
      end
    end
    if (reset) begin // @[ICache.scala 53:26]
      tag2_25 <= 53'h0; // @[ICache.scala 53:26]
    end else if (5'h19 == index_addr) begin // @[ICache.scala 99:26]
      if (_block2_T) begin // @[ICache.scala 99:32]
        tag2_25 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 57:28]
        tag2_25 <= tag2_31; // @[ICache.scala 57:28]
      end else begin
        tag2_25 <= _GEN_94;
      end
    end
    if (reset) begin // @[ICache.scala 53:26]
      tag2_26 <= 53'h0; // @[ICache.scala 53:26]
    end else if (5'h1a == index_addr) begin // @[ICache.scala 99:26]
      if (_block2_T) begin // @[ICache.scala 99:32]
        tag2_26 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 57:28]
        tag2_26 <= tag2_31; // @[ICache.scala 57:28]
      end else begin
        tag2_26 <= _GEN_94;
      end
    end
    if (reset) begin // @[ICache.scala 53:26]
      tag2_27 <= 53'h0; // @[ICache.scala 53:26]
    end else if (5'h1b == index_addr) begin // @[ICache.scala 99:26]
      if (_block2_T) begin // @[ICache.scala 99:32]
        tag2_27 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 57:28]
        tag2_27 <= tag2_31; // @[ICache.scala 57:28]
      end else begin
        tag2_27 <= _GEN_94;
      end
    end
    if (reset) begin // @[ICache.scala 53:26]
      tag2_28 <= 53'h0; // @[ICache.scala 53:26]
    end else if (5'h1c == index_addr) begin // @[ICache.scala 99:26]
      if (_block2_T) begin // @[ICache.scala 99:32]
        tag2_28 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 57:28]
        tag2_28 <= tag2_31; // @[ICache.scala 57:28]
      end else begin
        tag2_28 <= _GEN_94;
      end
    end
    if (reset) begin // @[ICache.scala 53:26]
      tag2_29 <= 53'h0; // @[ICache.scala 53:26]
    end else if (5'h1d == index_addr) begin // @[ICache.scala 99:26]
      if (_block2_T) begin // @[ICache.scala 99:32]
        tag2_29 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 57:28]
        tag2_29 <= tag2_31; // @[ICache.scala 57:28]
      end else begin
        tag2_29 <= _GEN_94;
      end
    end
    if (reset) begin // @[ICache.scala 53:26]
      tag2_30 <= 53'h0; // @[ICache.scala 53:26]
    end else if (5'h1e == index_addr) begin // @[ICache.scala 99:26]
      if (_block2_T) begin // @[ICache.scala 99:32]
        tag2_30 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 57:28]
        tag2_30 <= tag2_31; // @[ICache.scala 57:28]
      end else begin
        tag2_30 <= _GEN_94;
      end
    end
    if (reset) begin // @[ICache.scala 53:26]
      tag2_31 <= 53'h0; // @[ICache.scala 53:26]
    end else if (5'h1f == index_addr) begin // @[ICache.scala 99:26]
      if (_block2_T) begin // @[ICache.scala 99:32]
        tag2_31 <= tag_addr;
      end else if (!(5'h1f == index_addr)) begin // @[ICache.scala 57:28]
        tag2_31 <= _GEN_94;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      block2_0 <= 512'h0; // @[ICache.scala 54:26]
    end else if (5'h0 == index_addr) begin // @[ICache.scala 98:26]
      if (update & updateway2) begin // @[ICache.scala 98:32]
        block2_0 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 59:39]
        block2_0 <= block2_31; // @[ICache.scala 59:39]
      end else begin
        block2_0 <= _GEN_190;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      block2_1 <= 512'h0; // @[ICache.scala 54:26]
    end else if (5'h1 == index_addr) begin // @[ICache.scala 98:26]
      if (update & updateway2) begin // @[ICache.scala 98:32]
        block2_1 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 59:39]
        block2_1 <= block2_31; // @[ICache.scala 59:39]
      end else begin
        block2_1 <= _GEN_190;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      block2_2 <= 512'h0; // @[ICache.scala 54:26]
    end else if (5'h2 == index_addr) begin // @[ICache.scala 98:26]
      if (update & updateway2) begin // @[ICache.scala 98:32]
        block2_2 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 59:39]
        block2_2 <= block2_31; // @[ICache.scala 59:39]
      end else begin
        block2_2 <= _GEN_190;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      block2_3 <= 512'h0; // @[ICache.scala 54:26]
    end else if (5'h3 == index_addr) begin // @[ICache.scala 98:26]
      if (update & updateway2) begin // @[ICache.scala 98:32]
        block2_3 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 59:39]
        block2_3 <= block2_31; // @[ICache.scala 59:39]
      end else begin
        block2_3 <= _GEN_190;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      block2_4 <= 512'h0; // @[ICache.scala 54:26]
    end else if (5'h4 == index_addr) begin // @[ICache.scala 98:26]
      if (update & updateway2) begin // @[ICache.scala 98:32]
        block2_4 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 59:39]
        block2_4 <= block2_31; // @[ICache.scala 59:39]
      end else begin
        block2_4 <= _GEN_190;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      block2_5 <= 512'h0; // @[ICache.scala 54:26]
    end else if (5'h5 == index_addr) begin // @[ICache.scala 98:26]
      if (update & updateway2) begin // @[ICache.scala 98:32]
        block2_5 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 59:39]
        block2_5 <= block2_31; // @[ICache.scala 59:39]
      end else begin
        block2_5 <= _GEN_190;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      block2_6 <= 512'h0; // @[ICache.scala 54:26]
    end else if (5'h6 == index_addr) begin // @[ICache.scala 98:26]
      if (update & updateway2) begin // @[ICache.scala 98:32]
        block2_6 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 59:39]
        block2_6 <= block2_31; // @[ICache.scala 59:39]
      end else begin
        block2_6 <= _GEN_190;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      block2_7 <= 512'h0; // @[ICache.scala 54:26]
    end else if (5'h7 == index_addr) begin // @[ICache.scala 98:26]
      if (update & updateway2) begin // @[ICache.scala 98:32]
        block2_7 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 59:39]
        block2_7 <= block2_31; // @[ICache.scala 59:39]
      end else begin
        block2_7 <= _GEN_190;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      block2_8 <= 512'h0; // @[ICache.scala 54:26]
    end else if (5'h8 == index_addr) begin // @[ICache.scala 98:26]
      if (update & updateway2) begin // @[ICache.scala 98:32]
        block2_8 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 59:39]
        block2_8 <= block2_31; // @[ICache.scala 59:39]
      end else begin
        block2_8 <= _GEN_190;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      block2_9 <= 512'h0; // @[ICache.scala 54:26]
    end else if (5'h9 == index_addr) begin // @[ICache.scala 98:26]
      if (update & updateway2) begin // @[ICache.scala 98:32]
        block2_9 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 59:39]
        block2_9 <= block2_31; // @[ICache.scala 59:39]
      end else begin
        block2_9 <= _GEN_190;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      block2_10 <= 512'h0; // @[ICache.scala 54:26]
    end else if (5'ha == index_addr) begin // @[ICache.scala 98:26]
      if (update & updateway2) begin // @[ICache.scala 98:32]
        block2_10 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 59:39]
        block2_10 <= block2_31; // @[ICache.scala 59:39]
      end else begin
        block2_10 <= _GEN_190;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      block2_11 <= 512'h0; // @[ICache.scala 54:26]
    end else if (5'hb == index_addr) begin // @[ICache.scala 98:26]
      if (update & updateway2) begin // @[ICache.scala 98:32]
        block2_11 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 59:39]
        block2_11 <= block2_31; // @[ICache.scala 59:39]
      end else begin
        block2_11 <= _GEN_190;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      block2_12 <= 512'h0; // @[ICache.scala 54:26]
    end else if (5'hc == index_addr) begin // @[ICache.scala 98:26]
      if (update & updateway2) begin // @[ICache.scala 98:32]
        block2_12 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 59:39]
        block2_12 <= block2_31; // @[ICache.scala 59:39]
      end else begin
        block2_12 <= _GEN_190;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      block2_13 <= 512'h0; // @[ICache.scala 54:26]
    end else if (5'hd == index_addr) begin // @[ICache.scala 98:26]
      if (update & updateway2) begin // @[ICache.scala 98:32]
        block2_13 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 59:39]
        block2_13 <= block2_31; // @[ICache.scala 59:39]
      end else begin
        block2_13 <= _GEN_190;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      block2_14 <= 512'h0; // @[ICache.scala 54:26]
    end else if (5'he == index_addr) begin // @[ICache.scala 98:26]
      if (update & updateway2) begin // @[ICache.scala 98:32]
        block2_14 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 59:39]
        block2_14 <= block2_31; // @[ICache.scala 59:39]
      end else begin
        block2_14 <= _GEN_190;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      block2_15 <= 512'h0; // @[ICache.scala 54:26]
    end else if (5'hf == index_addr) begin // @[ICache.scala 98:26]
      if (update & updateway2) begin // @[ICache.scala 98:32]
        block2_15 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 59:39]
        block2_15 <= block2_31; // @[ICache.scala 59:39]
      end else begin
        block2_15 <= _GEN_190;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      block2_16 <= 512'h0; // @[ICache.scala 54:26]
    end else if (5'h10 == index_addr) begin // @[ICache.scala 98:26]
      if (update & updateway2) begin // @[ICache.scala 98:32]
        block2_16 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 59:39]
        block2_16 <= block2_31; // @[ICache.scala 59:39]
      end else begin
        block2_16 <= _GEN_190;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      block2_17 <= 512'h0; // @[ICache.scala 54:26]
    end else if (5'h11 == index_addr) begin // @[ICache.scala 98:26]
      if (update & updateway2) begin // @[ICache.scala 98:32]
        block2_17 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 59:39]
        block2_17 <= block2_31; // @[ICache.scala 59:39]
      end else begin
        block2_17 <= _GEN_190;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      block2_18 <= 512'h0; // @[ICache.scala 54:26]
    end else if (5'h12 == index_addr) begin // @[ICache.scala 98:26]
      if (update & updateway2) begin // @[ICache.scala 98:32]
        block2_18 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 59:39]
        block2_18 <= block2_31; // @[ICache.scala 59:39]
      end else begin
        block2_18 <= _GEN_190;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      block2_19 <= 512'h0; // @[ICache.scala 54:26]
    end else if (5'h13 == index_addr) begin // @[ICache.scala 98:26]
      if (update & updateway2) begin // @[ICache.scala 98:32]
        block2_19 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 59:39]
        block2_19 <= block2_31; // @[ICache.scala 59:39]
      end else begin
        block2_19 <= _GEN_190;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      block2_20 <= 512'h0; // @[ICache.scala 54:26]
    end else if (5'h14 == index_addr) begin // @[ICache.scala 98:26]
      if (update & updateway2) begin // @[ICache.scala 98:32]
        block2_20 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 59:39]
        block2_20 <= block2_31; // @[ICache.scala 59:39]
      end else begin
        block2_20 <= _GEN_190;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      block2_21 <= 512'h0; // @[ICache.scala 54:26]
    end else if (5'h15 == index_addr) begin // @[ICache.scala 98:26]
      if (update & updateway2) begin // @[ICache.scala 98:32]
        block2_21 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 59:39]
        block2_21 <= block2_31; // @[ICache.scala 59:39]
      end else begin
        block2_21 <= _GEN_190;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      block2_22 <= 512'h0; // @[ICache.scala 54:26]
    end else if (5'h16 == index_addr) begin // @[ICache.scala 98:26]
      if (update & updateway2) begin // @[ICache.scala 98:32]
        block2_22 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 59:39]
        block2_22 <= block2_31; // @[ICache.scala 59:39]
      end else begin
        block2_22 <= _GEN_190;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      block2_23 <= 512'h0; // @[ICache.scala 54:26]
    end else if (5'h17 == index_addr) begin // @[ICache.scala 98:26]
      if (update & updateway2) begin // @[ICache.scala 98:32]
        block2_23 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 59:39]
        block2_23 <= block2_31; // @[ICache.scala 59:39]
      end else begin
        block2_23 <= _GEN_190;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      block2_24 <= 512'h0; // @[ICache.scala 54:26]
    end else if (5'h18 == index_addr) begin // @[ICache.scala 98:26]
      if (update & updateway2) begin // @[ICache.scala 98:32]
        block2_24 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 59:39]
        block2_24 <= block2_31; // @[ICache.scala 59:39]
      end else begin
        block2_24 <= _GEN_190;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      block2_25 <= 512'h0; // @[ICache.scala 54:26]
    end else if (5'h19 == index_addr) begin // @[ICache.scala 98:26]
      if (update & updateway2) begin // @[ICache.scala 98:32]
        block2_25 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 59:39]
        block2_25 <= block2_31; // @[ICache.scala 59:39]
      end else begin
        block2_25 <= _GEN_190;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      block2_26 <= 512'h0; // @[ICache.scala 54:26]
    end else if (5'h1a == index_addr) begin // @[ICache.scala 98:26]
      if (update & updateway2) begin // @[ICache.scala 98:32]
        block2_26 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 59:39]
        block2_26 <= block2_31; // @[ICache.scala 59:39]
      end else begin
        block2_26 <= _GEN_190;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      block2_27 <= 512'h0; // @[ICache.scala 54:26]
    end else if (5'h1b == index_addr) begin // @[ICache.scala 98:26]
      if (update & updateway2) begin // @[ICache.scala 98:32]
        block2_27 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 59:39]
        block2_27 <= block2_31; // @[ICache.scala 59:39]
      end else begin
        block2_27 <= _GEN_190;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      block2_28 <= 512'h0; // @[ICache.scala 54:26]
    end else if (5'h1c == index_addr) begin // @[ICache.scala 98:26]
      if (update & updateway2) begin // @[ICache.scala 98:32]
        block2_28 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 59:39]
        block2_28 <= block2_31; // @[ICache.scala 59:39]
      end else begin
        block2_28 <= _GEN_190;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      block2_29 <= 512'h0; // @[ICache.scala 54:26]
    end else if (5'h1d == index_addr) begin // @[ICache.scala 98:26]
      if (update & updateway2) begin // @[ICache.scala 98:32]
        block2_29 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 59:39]
        block2_29 <= block2_31; // @[ICache.scala 59:39]
      end else begin
        block2_29 <= _GEN_190;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      block2_30 <= 512'h0; // @[ICache.scala 54:26]
    end else if (5'h1e == index_addr) begin // @[ICache.scala 98:26]
      if (update & updateway2) begin // @[ICache.scala 98:32]
        block2_30 <= io_axi_data;
      end else if (5'h1f == index_addr) begin // @[ICache.scala 59:39]
        block2_30 <= block2_31; // @[ICache.scala 59:39]
      end else begin
        block2_30 <= _GEN_190;
      end
    end
    if (reset) begin // @[ICache.scala 54:26]
      block2_31 <= 512'h0; // @[ICache.scala 54:26]
    end else if (5'h1f == index_addr) begin // @[ICache.scala 98:26]
      if (update & updateway2) begin // @[ICache.scala 98:32]
        block2_31 <= io_axi_data;
      end else if (!(5'h1f == index_addr)) begin // @[ICache.scala 59:39]
        block2_31 <= _GEN_190;
      end
    end
    if (hit2) begin // @[ICache.scala 62:22]
      io_imem_data_REG <= data2;
    end else if (hit1) begin // @[ICache.scala 62:39]
      io_imem_data_REG <= data1;
    end else begin
      io_imem_data_REG <= 32'h0;
    end
    io_imem_data_ok_REG <= reset | hit; // @[ICache.scala 70:31 ICache.scala 70:31 ICache.scala 70:31]
    if (reset) begin // @[ICache.scala 75:24]
      state <= 1'h0; // @[ICache.scala 75:24]
    end else if (_T) begin // @[Conditional.scala 40:58]
      state <= _GEN_320;
    end else if (state) begin // @[Conditional.scala 39:67]
      if (io_axi_valid) begin // @[ICache.scala 82:32]
        state <= 1'h0; // @[ICache.scala 82:39]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  v1_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  v1_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  v1_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  v1_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  v1_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  v1_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  v1_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  v1_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  v1_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  v1_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  v1_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  v1_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  v1_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  v1_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  v1_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  v1_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  v1_16 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  v1_17 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  v1_18 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  v1_19 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  v1_20 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  v1_21 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  v1_22 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  v1_23 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  v1_24 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  v1_25 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  v1_26 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  v1_27 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  v1_28 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  v1_29 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  v1_30 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  v1_31 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  age1_0 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  age1_1 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  age1_2 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  age1_3 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  age1_4 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  age1_5 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  age1_6 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  age1_7 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  age1_8 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  age1_9 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  age1_10 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  age1_11 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  age1_12 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  age1_13 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  age1_14 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  age1_15 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  age1_16 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  age1_17 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  age1_18 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  age1_19 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  age1_20 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  age1_21 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  age1_22 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  age1_23 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  age1_24 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  age1_25 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  age1_26 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  age1_27 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  age1_28 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  age1_29 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  age1_30 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  age1_31 = _RAND_63[0:0];
  _RAND_64 = {2{`RANDOM}};
  tag1_0 = _RAND_64[52:0];
  _RAND_65 = {2{`RANDOM}};
  tag1_1 = _RAND_65[52:0];
  _RAND_66 = {2{`RANDOM}};
  tag1_2 = _RAND_66[52:0];
  _RAND_67 = {2{`RANDOM}};
  tag1_3 = _RAND_67[52:0];
  _RAND_68 = {2{`RANDOM}};
  tag1_4 = _RAND_68[52:0];
  _RAND_69 = {2{`RANDOM}};
  tag1_5 = _RAND_69[52:0];
  _RAND_70 = {2{`RANDOM}};
  tag1_6 = _RAND_70[52:0];
  _RAND_71 = {2{`RANDOM}};
  tag1_7 = _RAND_71[52:0];
  _RAND_72 = {2{`RANDOM}};
  tag1_8 = _RAND_72[52:0];
  _RAND_73 = {2{`RANDOM}};
  tag1_9 = _RAND_73[52:0];
  _RAND_74 = {2{`RANDOM}};
  tag1_10 = _RAND_74[52:0];
  _RAND_75 = {2{`RANDOM}};
  tag1_11 = _RAND_75[52:0];
  _RAND_76 = {2{`RANDOM}};
  tag1_12 = _RAND_76[52:0];
  _RAND_77 = {2{`RANDOM}};
  tag1_13 = _RAND_77[52:0];
  _RAND_78 = {2{`RANDOM}};
  tag1_14 = _RAND_78[52:0];
  _RAND_79 = {2{`RANDOM}};
  tag1_15 = _RAND_79[52:0];
  _RAND_80 = {2{`RANDOM}};
  tag1_16 = _RAND_80[52:0];
  _RAND_81 = {2{`RANDOM}};
  tag1_17 = _RAND_81[52:0];
  _RAND_82 = {2{`RANDOM}};
  tag1_18 = _RAND_82[52:0];
  _RAND_83 = {2{`RANDOM}};
  tag1_19 = _RAND_83[52:0];
  _RAND_84 = {2{`RANDOM}};
  tag1_20 = _RAND_84[52:0];
  _RAND_85 = {2{`RANDOM}};
  tag1_21 = _RAND_85[52:0];
  _RAND_86 = {2{`RANDOM}};
  tag1_22 = _RAND_86[52:0];
  _RAND_87 = {2{`RANDOM}};
  tag1_23 = _RAND_87[52:0];
  _RAND_88 = {2{`RANDOM}};
  tag1_24 = _RAND_88[52:0];
  _RAND_89 = {2{`RANDOM}};
  tag1_25 = _RAND_89[52:0];
  _RAND_90 = {2{`RANDOM}};
  tag1_26 = _RAND_90[52:0];
  _RAND_91 = {2{`RANDOM}};
  tag1_27 = _RAND_91[52:0];
  _RAND_92 = {2{`RANDOM}};
  tag1_28 = _RAND_92[52:0];
  _RAND_93 = {2{`RANDOM}};
  tag1_29 = _RAND_93[52:0];
  _RAND_94 = {2{`RANDOM}};
  tag1_30 = _RAND_94[52:0];
  _RAND_95 = {2{`RANDOM}};
  tag1_31 = _RAND_95[52:0];
  _RAND_96 = {16{`RANDOM}};
  block1_0 = _RAND_96[511:0];
  _RAND_97 = {16{`RANDOM}};
  block1_1 = _RAND_97[511:0];
  _RAND_98 = {16{`RANDOM}};
  block1_2 = _RAND_98[511:0];
  _RAND_99 = {16{`RANDOM}};
  block1_3 = _RAND_99[511:0];
  _RAND_100 = {16{`RANDOM}};
  block1_4 = _RAND_100[511:0];
  _RAND_101 = {16{`RANDOM}};
  block1_5 = _RAND_101[511:0];
  _RAND_102 = {16{`RANDOM}};
  block1_6 = _RAND_102[511:0];
  _RAND_103 = {16{`RANDOM}};
  block1_7 = _RAND_103[511:0];
  _RAND_104 = {16{`RANDOM}};
  block1_8 = _RAND_104[511:0];
  _RAND_105 = {16{`RANDOM}};
  block1_9 = _RAND_105[511:0];
  _RAND_106 = {16{`RANDOM}};
  block1_10 = _RAND_106[511:0];
  _RAND_107 = {16{`RANDOM}};
  block1_11 = _RAND_107[511:0];
  _RAND_108 = {16{`RANDOM}};
  block1_12 = _RAND_108[511:0];
  _RAND_109 = {16{`RANDOM}};
  block1_13 = _RAND_109[511:0];
  _RAND_110 = {16{`RANDOM}};
  block1_14 = _RAND_110[511:0];
  _RAND_111 = {16{`RANDOM}};
  block1_15 = _RAND_111[511:0];
  _RAND_112 = {16{`RANDOM}};
  block1_16 = _RAND_112[511:0];
  _RAND_113 = {16{`RANDOM}};
  block1_17 = _RAND_113[511:0];
  _RAND_114 = {16{`RANDOM}};
  block1_18 = _RAND_114[511:0];
  _RAND_115 = {16{`RANDOM}};
  block1_19 = _RAND_115[511:0];
  _RAND_116 = {16{`RANDOM}};
  block1_20 = _RAND_116[511:0];
  _RAND_117 = {16{`RANDOM}};
  block1_21 = _RAND_117[511:0];
  _RAND_118 = {16{`RANDOM}};
  block1_22 = _RAND_118[511:0];
  _RAND_119 = {16{`RANDOM}};
  block1_23 = _RAND_119[511:0];
  _RAND_120 = {16{`RANDOM}};
  block1_24 = _RAND_120[511:0];
  _RAND_121 = {16{`RANDOM}};
  block1_25 = _RAND_121[511:0];
  _RAND_122 = {16{`RANDOM}};
  block1_26 = _RAND_122[511:0];
  _RAND_123 = {16{`RANDOM}};
  block1_27 = _RAND_123[511:0];
  _RAND_124 = {16{`RANDOM}};
  block1_28 = _RAND_124[511:0];
  _RAND_125 = {16{`RANDOM}};
  block1_29 = _RAND_125[511:0];
  _RAND_126 = {16{`RANDOM}};
  block1_30 = _RAND_126[511:0];
  _RAND_127 = {16{`RANDOM}};
  block1_31 = _RAND_127[511:0];
  _RAND_128 = {1{`RANDOM}};
  v2_0 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  v2_1 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  v2_2 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  v2_3 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  v2_4 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  v2_5 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  v2_6 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  v2_7 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  v2_8 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  v2_9 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  v2_10 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  v2_11 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  v2_12 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  v2_13 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  v2_14 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  v2_15 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  v2_16 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  v2_17 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  v2_18 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  v2_19 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  v2_20 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  v2_21 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  v2_22 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  v2_23 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  v2_24 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  v2_25 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  v2_26 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  v2_27 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  v2_28 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  v2_29 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  v2_30 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  v2_31 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  age2_0 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  age2_1 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  age2_2 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  age2_3 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  age2_4 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  age2_5 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  age2_6 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  age2_7 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  age2_8 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  age2_9 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  age2_10 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  age2_11 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  age2_12 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  age2_13 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  age2_14 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  age2_15 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  age2_16 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  age2_17 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  age2_18 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  age2_19 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  age2_20 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  age2_21 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  age2_22 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  age2_23 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  age2_24 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  age2_25 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  age2_26 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  age2_27 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  age2_28 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  age2_29 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  age2_30 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  age2_31 = _RAND_191[0:0];
  _RAND_192 = {2{`RANDOM}};
  tag2_0 = _RAND_192[52:0];
  _RAND_193 = {2{`RANDOM}};
  tag2_1 = _RAND_193[52:0];
  _RAND_194 = {2{`RANDOM}};
  tag2_2 = _RAND_194[52:0];
  _RAND_195 = {2{`RANDOM}};
  tag2_3 = _RAND_195[52:0];
  _RAND_196 = {2{`RANDOM}};
  tag2_4 = _RAND_196[52:0];
  _RAND_197 = {2{`RANDOM}};
  tag2_5 = _RAND_197[52:0];
  _RAND_198 = {2{`RANDOM}};
  tag2_6 = _RAND_198[52:0];
  _RAND_199 = {2{`RANDOM}};
  tag2_7 = _RAND_199[52:0];
  _RAND_200 = {2{`RANDOM}};
  tag2_8 = _RAND_200[52:0];
  _RAND_201 = {2{`RANDOM}};
  tag2_9 = _RAND_201[52:0];
  _RAND_202 = {2{`RANDOM}};
  tag2_10 = _RAND_202[52:0];
  _RAND_203 = {2{`RANDOM}};
  tag2_11 = _RAND_203[52:0];
  _RAND_204 = {2{`RANDOM}};
  tag2_12 = _RAND_204[52:0];
  _RAND_205 = {2{`RANDOM}};
  tag2_13 = _RAND_205[52:0];
  _RAND_206 = {2{`RANDOM}};
  tag2_14 = _RAND_206[52:0];
  _RAND_207 = {2{`RANDOM}};
  tag2_15 = _RAND_207[52:0];
  _RAND_208 = {2{`RANDOM}};
  tag2_16 = _RAND_208[52:0];
  _RAND_209 = {2{`RANDOM}};
  tag2_17 = _RAND_209[52:0];
  _RAND_210 = {2{`RANDOM}};
  tag2_18 = _RAND_210[52:0];
  _RAND_211 = {2{`RANDOM}};
  tag2_19 = _RAND_211[52:0];
  _RAND_212 = {2{`RANDOM}};
  tag2_20 = _RAND_212[52:0];
  _RAND_213 = {2{`RANDOM}};
  tag2_21 = _RAND_213[52:0];
  _RAND_214 = {2{`RANDOM}};
  tag2_22 = _RAND_214[52:0];
  _RAND_215 = {2{`RANDOM}};
  tag2_23 = _RAND_215[52:0];
  _RAND_216 = {2{`RANDOM}};
  tag2_24 = _RAND_216[52:0];
  _RAND_217 = {2{`RANDOM}};
  tag2_25 = _RAND_217[52:0];
  _RAND_218 = {2{`RANDOM}};
  tag2_26 = _RAND_218[52:0];
  _RAND_219 = {2{`RANDOM}};
  tag2_27 = _RAND_219[52:0];
  _RAND_220 = {2{`RANDOM}};
  tag2_28 = _RAND_220[52:0];
  _RAND_221 = {2{`RANDOM}};
  tag2_29 = _RAND_221[52:0];
  _RAND_222 = {2{`RANDOM}};
  tag2_30 = _RAND_222[52:0];
  _RAND_223 = {2{`RANDOM}};
  tag2_31 = _RAND_223[52:0];
  _RAND_224 = {16{`RANDOM}};
  block2_0 = _RAND_224[511:0];
  _RAND_225 = {16{`RANDOM}};
  block2_1 = _RAND_225[511:0];
  _RAND_226 = {16{`RANDOM}};
  block2_2 = _RAND_226[511:0];
  _RAND_227 = {16{`RANDOM}};
  block2_3 = _RAND_227[511:0];
  _RAND_228 = {16{`RANDOM}};
  block2_4 = _RAND_228[511:0];
  _RAND_229 = {16{`RANDOM}};
  block2_5 = _RAND_229[511:0];
  _RAND_230 = {16{`RANDOM}};
  block2_6 = _RAND_230[511:0];
  _RAND_231 = {16{`RANDOM}};
  block2_7 = _RAND_231[511:0];
  _RAND_232 = {16{`RANDOM}};
  block2_8 = _RAND_232[511:0];
  _RAND_233 = {16{`RANDOM}};
  block2_9 = _RAND_233[511:0];
  _RAND_234 = {16{`RANDOM}};
  block2_10 = _RAND_234[511:0];
  _RAND_235 = {16{`RANDOM}};
  block2_11 = _RAND_235[511:0];
  _RAND_236 = {16{`RANDOM}};
  block2_12 = _RAND_236[511:0];
  _RAND_237 = {16{`RANDOM}};
  block2_13 = _RAND_237[511:0];
  _RAND_238 = {16{`RANDOM}};
  block2_14 = _RAND_238[511:0];
  _RAND_239 = {16{`RANDOM}};
  block2_15 = _RAND_239[511:0];
  _RAND_240 = {16{`RANDOM}};
  block2_16 = _RAND_240[511:0];
  _RAND_241 = {16{`RANDOM}};
  block2_17 = _RAND_241[511:0];
  _RAND_242 = {16{`RANDOM}};
  block2_18 = _RAND_242[511:0];
  _RAND_243 = {16{`RANDOM}};
  block2_19 = _RAND_243[511:0];
  _RAND_244 = {16{`RANDOM}};
  block2_20 = _RAND_244[511:0];
  _RAND_245 = {16{`RANDOM}};
  block2_21 = _RAND_245[511:0];
  _RAND_246 = {16{`RANDOM}};
  block2_22 = _RAND_246[511:0];
  _RAND_247 = {16{`RANDOM}};
  block2_23 = _RAND_247[511:0];
  _RAND_248 = {16{`RANDOM}};
  block2_24 = _RAND_248[511:0];
  _RAND_249 = {16{`RANDOM}};
  block2_25 = _RAND_249[511:0];
  _RAND_250 = {16{`RANDOM}};
  block2_26 = _RAND_250[511:0];
  _RAND_251 = {16{`RANDOM}};
  block2_27 = _RAND_251[511:0];
  _RAND_252 = {16{`RANDOM}};
  block2_28 = _RAND_252[511:0];
  _RAND_253 = {16{`RANDOM}};
  block2_29 = _RAND_253[511:0];
  _RAND_254 = {16{`RANDOM}};
  block2_30 = _RAND_254[511:0];
  _RAND_255 = {16{`RANDOM}};
  block2_31 = _RAND_255[511:0];
  _RAND_256 = {1{`RANDOM}};
  io_imem_data_REG = _RAND_256[31:0];
  _RAND_257 = {1{`RANDOM}};
  io_imem_data_ok_REG = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  state = _RAND_258[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DCache(
  input          clock,
  input          reset,
  input          io_dmem_en,
  input          io_dmem_op,
  input  [63:0]  io_dmem_addr,
  input  [63:0]  io_dmem_wdata,
  input  [7:0]   io_dmem_wmask,
  output         io_dmem_ok,
  output [63:0]  io_dmem_rdata,
  output         io_axi_req,
  output [63:0]  io_axi_raddr,
  input          io_axi_rvalid,
  input  [511:0] io_axi_rdata,
  output         io_axi_weq,
  output [63:0]  io_axi_waddr,
  output [511:0] io_axi_wdata,
  input          io_axi_wdone
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [63:0] _RAND_100;
  reg [63:0] _RAND_101;
  reg [63:0] _RAND_102;
  reg [63:0] _RAND_103;
  reg [63:0] _RAND_104;
  reg [63:0] _RAND_105;
  reg [63:0] _RAND_106;
  reg [63:0] _RAND_107;
  reg [63:0] _RAND_108;
  reg [63:0] _RAND_109;
  reg [63:0] _RAND_110;
  reg [63:0] _RAND_111;
  reg [63:0] _RAND_112;
  reg [63:0] _RAND_113;
  reg [63:0] _RAND_114;
  reg [63:0] _RAND_115;
  reg [63:0] _RAND_116;
  reg [63:0] _RAND_117;
  reg [63:0] _RAND_118;
  reg [63:0] _RAND_119;
  reg [63:0] _RAND_120;
  reg [63:0] _RAND_121;
  reg [63:0] _RAND_122;
  reg [63:0] _RAND_123;
  reg [63:0] _RAND_124;
  reg [63:0] _RAND_125;
  reg [63:0] _RAND_126;
  reg [63:0] _RAND_127;
  reg [63:0] _RAND_128;
  reg [63:0] _RAND_129;
  reg [63:0] _RAND_130;
  reg [63:0] _RAND_131;
  reg [511:0] _RAND_132;
  reg [511:0] _RAND_133;
  reg [511:0] _RAND_134;
  reg [511:0] _RAND_135;
  reg [511:0] _RAND_136;
  reg [511:0] _RAND_137;
  reg [511:0] _RAND_138;
  reg [511:0] _RAND_139;
  reg [511:0] _RAND_140;
  reg [511:0] _RAND_141;
  reg [511:0] _RAND_142;
  reg [511:0] _RAND_143;
  reg [511:0] _RAND_144;
  reg [511:0] _RAND_145;
  reg [511:0] _RAND_146;
  reg [511:0] _RAND_147;
  reg [511:0] _RAND_148;
  reg [511:0] _RAND_149;
  reg [511:0] _RAND_150;
  reg [511:0] _RAND_151;
  reg [511:0] _RAND_152;
  reg [511:0] _RAND_153;
  reg [511:0] _RAND_154;
  reg [511:0] _RAND_155;
  reg [511:0] _RAND_156;
  reg [511:0] _RAND_157;
  reg [511:0] _RAND_158;
  reg [511:0] _RAND_159;
  reg [511:0] _RAND_160;
  reg [511:0] _RAND_161;
  reg [511:0] _RAND_162;
  reg [511:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [63:0] _RAND_260;
  reg [63:0] _RAND_261;
  reg [63:0] _RAND_262;
  reg [63:0] _RAND_263;
  reg [63:0] _RAND_264;
  reg [63:0] _RAND_265;
  reg [63:0] _RAND_266;
  reg [63:0] _RAND_267;
  reg [63:0] _RAND_268;
  reg [63:0] _RAND_269;
  reg [63:0] _RAND_270;
  reg [63:0] _RAND_271;
  reg [63:0] _RAND_272;
  reg [63:0] _RAND_273;
  reg [63:0] _RAND_274;
  reg [63:0] _RAND_275;
  reg [63:0] _RAND_276;
  reg [63:0] _RAND_277;
  reg [63:0] _RAND_278;
  reg [63:0] _RAND_279;
  reg [63:0] _RAND_280;
  reg [63:0] _RAND_281;
  reg [63:0] _RAND_282;
  reg [63:0] _RAND_283;
  reg [63:0] _RAND_284;
  reg [63:0] _RAND_285;
  reg [63:0] _RAND_286;
  reg [63:0] _RAND_287;
  reg [63:0] _RAND_288;
  reg [63:0] _RAND_289;
  reg [63:0] _RAND_290;
  reg [63:0] _RAND_291;
  reg [511:0] _RAND_292;
  reg [511:0] _RAND_293;
  reg [511:0] _RAND_294;
  reg [511:0] _RAND_295;
  reg [511:0] _RAND_296;
  reg [511:0] _RAND_297;
  reg [511:0] _RAND_298;
  reg [511:0] _RAND_299;
  reg [511:0] _RAND_300;
  reg [511:0] _RAND_301;
  reg [511:0] _RAND_302;
  reg [511:0] _RAND_303;
  reg [511:0] _RAND_304;
  reg [511:0] _RAND_305;
  reg [511:0] _RAND_306;
  reg [511:0] _RAND_307;
  reg [511:0] _RAND_308;
  reg [511:0] _RAND_309;
  reg [511:0] _RAND_310;
  reg [511:0] _RAND_311;
  reg [511:0] _RAND_312;
  reg [511:0] _RAND_313;
  reg [511:0] _RAND_314;
  reg [511:0] _RAND_315;
  reg [511:0] _RAND_316;
  reg [511:0] _RAND_317;
  reg [511:0] _RAND_318;
  reg [511:0] _RAND_319;
  reg [511:0] _RAND_320;
  reg [511:0] _RAND_321;
  reg [511:0] _RAND_322;
  reg [511:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
`endif // RANDOMIZE_REG_INIT
  wire  _op_T = io_dmem_en & io_dmem_ok; // @[DCache.scala 39:66]
  reg  op; // @[Reg.scala 27:20]
  reg [63:0] addr; // @[Reg.scala 27:20]
  reg [63:0] wdata; // @[Reg.scala 27:20]
  reg [7:0] wm; // @[Reg.scala 27:20]
  wire [52:0] tag_addr = addr[63:11]; // @[DCache.scala 45:27]
  wire [4:0] index_addr = addr[10:6]; // @[DCache.scala 46:27]
  wire [5:0] offset_addr = addr[5:0]; // @[DCache.scala 47:27]
  reg  v1_0; // @[DCache.scala 49:26]
  reg  v1_1; // @[DCache.scala 49:26]
  reg  v1_2; // @[DCache.scala 49:26]
  reg  v1_3; // @[DCache.scala 49:26]
  reg  v1_4; // @[DCache.scala 49:26]
  reg  v1_5; // @[DCache.scala 49:26]
  reg  v1_6; // @[DCache.scala 49:26]
  reg  v1_7; // @[DCache.scala 49:26]
  reg  v1_8; // @[DCache.scala 49:26]
  reg  v1_9; // @[DCache.scala 49:26]
  reg  v1_10; // @[DCache.scala 49:26]
  reg  v1_11; // @[DCache.scala 49:26]
  reg  v1_12; // @[DCache.scala 49:26]
  reg  v1_13; // @[DCache.scala 49:26]
  reg  v1_14; // @[DCache.scala 49:26]
  reg  v1_15; // @[DCache.scala 49:26]
  reg  v1_16; // @[DCache.scala 49:26]
  reg  v1_17; // @[DCache.scala 49:26]
  reg  v1_18; // @[DCache.scala 49:26]
  reg  v1_19; // @[DCache.scala 49:26]
  reg  v1_20; // @[DCache.scala 49:26]
  reg  v1_21; // @[DCache.scala 49:26]
  reg  v1_22; // @[DCache.scala 49:26]
  reg  v1_23; // @[DCache.scala 49:26]
  reg  v1_24; // @[DCache.scala 49:26]
  reg  v1_25; // @[DCache.scala 49:26]
  reg  v1_26; // @[DCache.scala 49:26]
  reg  v1_27; // @[DCache.scala 49:26]
  reg  v1_28; // @[DCache.scala 49:26]
  reg  v1_29; // @[DCache.scala 49:26]
  reg  v1_30; // @[DCache.scala 49:26]
  reg  v1_31; // @[DCache.scala 49:26]
  reg  d1_0; // @[DCache.scala 50:26]
  reg  d1_1; // @[DCache.scala 50:26]
  reg  d1_2; // @[DCache.scala 50:26]
  reg  d1_3; // @[DCache.scala 50:26]
  reg  d1_4; // @[DCache.scala 50:26]
  reg  d1_5; // @[DCache.scala 50:26]
  reg  d1_6; // @[DCache.scala 50:26]
  reg  d1_7; // @[DCache.scala 50:26]
  reg  d1_8; // @[DCache.scala 50:26]
  reg  d1_9; // @[DCache.scala 50:26]
  reg  d1_10; // @[DCache.scala 50:26]
  reg  d1_11; // @[DCache.scala 50:26]
  reg  d1_12; // @[DCache.scala 50:26]
  reg  d1_13; // @[DCache.scala 50:26]
  reg  d1_14; // @[DCache.scala 50:26]
  reg  d1_15; // @[DCache.scala 50:26]
  reg  d1_16; // @[DCache.scala 50:26]
  reg  d1_17; // @[DCache.scala 50:26]
  reg  d1_18; // @[DCache.scala 50:26]
  reg  d1_19; // @[DCache.scala 50:26]
  reg  d1_20; // @[DCache.scala 50:26]
  reg  d1_21; // @[DCache.scala 50:26]
  reg  d1_22; // @[DCache.scala 50:26]
  reg  d1_23; // @[DCache.scala 50:26]
  reg  d1_24; // @[DCache.scala 50:26]
  reg  d1_25; // @[DCache.scala 50:26]
  reg  d1_26; // @[DCache.scala 50:26]
  reg  d1_27; // @[DCache.scala 50:26]
  reg  d1_28; // @[DCache.scala 50:26]
  reg  d1_29; // @[DCache.scala 50:26]
  reg  d1_30; // @[DCache.scala 50:26]
  reg  d1_31; // @[DCache.scala 50:26]
  reg  age1_0; // @[DCache.scala 51:26]
  reg  age1_1; // @[DCache.scala 51:26]
  reg  age1_2; // @[DCache.scala 51:26]
  reg  age1_3; // @[DCache.scala 51:26]
  reg  age1_4; // @[DCache.scala 51:26]
  reg  age1_5; // @[DCache.scala 51:26]
  reg  age1_6; // @[DCache.scala 51:26]
  reg  age1_7; // @[DCache.scala 51:26]
  reg  age1_8; // @[DCache.scala 51:26]
  reg  age1_9; // @[DCache.scala 51:26]
  reg  age1_10; // @[DCache.scala 51:26]
  reg  age1_11; // @[DCache.scala 51:26]
  reg  age1_12; // @[DCache.scala 51:26]
  reg  age1_13; // @[DCache.scala 51:26]
  reg  age1_14; // @[DCache.scala 51:26]
  reg  age1_15; // @[DCache.scala 51:26]
  reg  age1_16; // @[DCache.scala 51:26]
  reg  age1_17; // @[DCache.scala 51:26]
  reg  age1_18; // @[DCache.scala 51:26]
  reg  age1_19; // @[DCache.scala 51:26]
  reg  age1_20; // @[DCache.scala 51:26]
  reg  age1_21; // @[DCache.scala 51:26]
  reg  age1_22; // @[DCache.scala 51:26]
  reg  age1_23; // @[DCache.scala 51:26]
  reg  age1_24; // @[DCache.scala 51:26]
  reg  age1_25; // @[DCache.scala 51:26]
  reg  age1_26; // @[DCache.scala 51:26]
  reg  age1_27; // @[DCache.scala 51:26]
  reg  age1_28; // @[DCache.scala 51:26]
  reg  age1_29; // @[DCache.scala 51:26]
  reg  age1_30; // @[DCache.scala 51:26]
  reg  age1_31; // @[DCache.scala 51:26]
  reg [52:0] tag1_0; // @[DCache.scala 52:26]
  reg [52:0] tag1_1; // @[DCache.scala 52:26]
  reg [52:0] tag1_2; // @[DCache.scala 52:26]
  reg [52:0] tag1_3; // @[DCache.scala 52:26]
  reg [52:0] tag1_4; // @[DCache.scala 52:26]
  reg [52:0] tag1_5; // @[DCache.scala 52:26]
  reg [52:0] tag1_6; // @[DCache.scala 52:26]
  reg [52:0] tag1_7; // @[DCache.scala 52:26]
  reg [52:0] tag1_8; // @[DCache.scala 52:26]
  reg [52:0] tag1_9; // @[DCache.scala 52:26]
  reg [52:0] tag1_10; // @[DCache.scala 52:26]
  reg [52:0] tag1_11; // @[DCache.scala 52:26]
  reg [52:0] tag1_12; // @[DCache.scala 52:26]
  reg [52:0] tag1_13; // @[DCache.scala 52:26]
  reg [52:0] tag1_14; // @[DCache.scala 52:26]
  reg [52:0] tag1_15; // @[DCache.scala 52:26]
  reg [52:0] tag1_16; // @[DCache.scala 52:26]
  reg [52:0] tag1_17; // @[DCache.scala 52:26]
  reg [52:0] tag1_18; // @[DCache.scala 52:26]
  reg [52:0] tag1_19; // @[DCache.scala 52:26]
  reg [52:0] tag1_20; // @[DCache.scala 52:26]
  reg [52:0] tag1_21; // @[DCache.scala 52:26]
  reg [52:0] tag1_22; // @[DCache.scala 52:26]
  reg [52:0] tag1_23; // @[DCache.scala 52:26]
  reg [52:0] tag1_24; // @[DCache.scala 52:26]
  reg [52:0] tag1_25; // @[DCache.scala 52:26]
  reg [52:0] tag1_26; // @[DCache.scala 52:26]
  reg [52:0] tag1_27; // @[DCache.scala 52:26]
  reg [52:0] tag1_28; // @[DCache.scala 52:26]
  reg [52:0] tag1_29; // @[DCache.scala 52:26]
  reg [52:0] tag1_30; // @[DCache.scala 52:26]
  reg [52:0] tag1_31; // @[DCache.scala 52:26]
  reg [511:0] block1_0; // @[DCache.scala 53:26]
  reg [511:0] block1_1; // @[DCache.scala 53:26]
  reg [511:0] block1_2; // @[DCache.scala 53:26]
  reg [511:0] block1_3; // @[DCache.scala 53:26]
  reg [511:0] block1_4; // @[DCache.scala 53:26]
  reg [511:0] block1_5; // @[DCache.scala 53:26]
  reg [511:0] block1_6; // @[DCache.scala 53:26]
  reg [511:0] block1_7; // @[DCache.scala 53:26]
  reg [511:0] block1_8; // @[DCache.scala 53:26]
  reg [511:0] block1_9; // @[DCache.scala 53:26]
  reg [511:0] block1_10; // @[DCache.scala 53:26]
  reg [511:0] block1_11; // @[DCache.scala 53:26]
  reg [511:0] block1_12; // @[DCache.scala 53:26]
  reg [511:0] block1_13; // @[DCache.scala 53:26]
  reg [511:0] block1_14; // @[DCache.scala 53:26]
  reg [511:0] block1_15; // @[DCache.scala 53:26]
  reg [511:0] block1_16; // @[DCache.scala 53:26]
  reg [511:0] block1_17; // @[DCache.scala 53:26]
  reg [511:0] block1_18; // @[DCache.scala 53:26]
  reg [511:0] block1_19; // @[DCache.scala 53:26]
  reg [511:0] block1_20; // @[DCache.scala 53:26]
  reg [511:0] block1_21; // @[DCache.scala 53:26]
  reg [511:0] block1_22; // @[DCache.scala 53:26]
  reg [511:0] block1_23; // @[DCache.scala 53:26]
  reg [511:0] block1_24; // @[DCache.scala 53:26]
  reg [511:0] block1_25; // @[DCache.scala 53:26]
  reg [511:0] block1_26; // @[DCache.scala 53:26]
  reg [511:0] block1_27; // @[DCache.scala 53:26]
  reg [511:0] block1_28; // @[DCache.scala 53:26]
  reg [511:0] block1_29; // @[DCache.scala 53:26]
  reg [511:0] block1_30; // @[DCache.scala 53:26]
  reg [511:0] block1_31; // @[DCache.scala 53:26]
  reg  v2_0; // @[DCache.scala 54:26]
  reg  v2_1; // @[DCache.scala 54:26]
  reg  v2_2; // @[DCache.scala 54:26]
  reg  v2_3; // @[DCache.scala 54:26]
  reg  v2_4; // @[DCache.scala 54:26]
  reg  v2_5; // @[DCache.scala 54:26]
  reg  v2_6; // @[DCache.scala 54:26]
  reg  v2_7; // @[DCache.scala 54:26]
  reg  v2_8; // @[DCache.scala 54:26]
  reg  v2_9; // @[DCache.scala 54:26]
  reg  v2_10; // @[DCache.scala 54:26]
  reg  v2_11; // @[DCache.scala 54:26]
  reg  v2_12; // @[DCache.scala 54:26]
  reg  v2_13; // @[DCache.scala 54:26]
  reg  v2_14; // @[DCache.scala 54:26]
  reg  v2_15; // @[DCache.scala 54:26]
  reg  v2_16; // @[DCache.scala 54:26]
  reg  v2_17; // @[DCache.scala 54:26]
  reg  v2_18; // @[DCache.scala 54:26]
  reg  v2_19; // @[DCache.scala 54:26]
  reg  v2_20; // @[DCache.scala 54:26]
  reg  v2_21; // @[DCache.scala 54:26]
  reg  v2_22; // @[DCache.scala 54:26]
  reg  v2_23; // @[DCache.scala 54:26]
  reg  v2_24; // @[DCache.scala 54:26]
  reg  v2_25; // @[DCache.scala 54:26]
  reg  v2_26; // @[DCache.scala 54:26]
  reg  v2_27; // @[DCache.scala 54:26]
  reg  v2_28; // @[DCache.scala 54:26]
  reg  v2_29; // @[DCache.scala 54:26]
  reg  v2_30; // @[DCache.scala 54:26]
  reg  v2_31; // @[DCache.scala 54:26]
  reg  d2_0; // @[DCache.scala 55:26]
  reg  d2_1; // @[DCache.scala 55:26]
  reg  d2_2; // @[DCache.scala 55:26]
  reg  d2_3; // @[DCache.scala 55:26]
  reg  d2_4; // @[DCache.scala 55:26]
  reg  d2_5; // @[DCache.scala 55:26]
  reg  d2_6; // @[DCache.scala 55:26]
  reg  d2_7; // @[DCache.scala 55:26]
  reg  d2_8; // @[DCache.scala 55:26]
  reg  d2_9; // @[DCache.scala 55:26]
  reg  d2_10; // @[DCache.scala 55:26]
  reg  d2_11; // @[DCache.scala 55:26]
  reg  d2_12; // @[DCache.scala 55:26]
  reg  d2_13; // @[DCache.scala 55:26]
  reg  d2_14; // @[DCache.scala 55:26]
  reg  d2_15; // @[DCache.scala 55:26]
  reg  d2_16; // @[DCache.scala 55:26]
  reg  d2_17; // @[DCache.scala 55:26]
  reg  d2_18; // @[DCache.scala 55:26]
  reg  d2_19; // @[DCache.scala 55:26]
  reg  d2_20; // @[DCache.scala 55:26]
  reg  d2_21; // @[DCache.scala 55:26]
  reg  d2_22; // @[DCache.scala 55:26]
  reg  d2_23; // @[DCache.scala 55:26]
  reg  d2_24; // @[DCache.scala 55:26]
  reg  d2_25; // @[DCache.scala 55:26]
  reg  d2_26; // @[DCache.scala 55:26]
  reg  d2_27; // @[DCache.scala 55:26]
  reg  d2_28; // @[DCache.scala 55:26]
  reg  d2_29; // @[DCache.scala 55:26]
  reg  d2_30; // @[DCache.scala 55:26]
  reg  d2_31; // @[DCache.scala 55:26]
  reg  age2_0; // @[DCache.scala 56:26]
  reg  age2_1; // @[DCache.scala 56:26]
  reg  age2_2; // @[DCache.scala 56:26]
  reg  age2_3; // @[DCache.scala 56:26]
  reg  age2_4; // @[DCache.scala 56:26]
  reg  age2_5; // @[DCache.scala 56:26]
  reg  age2_6; // @[DCache.scala 56:26]
  reg  age2_7; // @[DCache.scala 56:26]
  reg  age2_8; // @[DCache.scala 56:26]
  reg  age2_9; // @[DCache.scala 56:26]
  reg  age2_10; // @[DCache.scala 56:26]
  reg  age2_11; // @[DCache.scala 56:26]
  reg  age2_12; // @[DCache.scala 56:26]
  reg  age2_13; // @[DCache.scala 56:26]
  reg  age2_14; // @[DCache.scala 56:26]
  reg  age2_15; // @[DCache.scala 56:26]
  reg  age2_16; // @[DCache.scala 56:26]
  reg  age2_17; // @[DCache.scala 56:26]
  reg  age2_18; // @[DCache.scala 56:26]
  reg  age2_19; // @[DCache.scala 56:26]
  reg  age2_20; // @[DCache.scala 56:26]
  reg  age2_21; // @[DCache.scala 56:26]
  reg  age2_22; // @[DCache.scala 56:26]
  reg  age2_23; // @[DCache.scala 56:26]
  reg  age2_24; // @[DCache.scala 56:26]
  reg  age2_25; // @[DCache.scala 56:26]
  reg  age2_26; // @[DCache.scala 56:26]
  reg  age2_27; // @[DCache.scala 56:26]
  reg  age2_28; // @[DCache.scala 56:26]
  reg  age2_29; // @[DCache.scala 56:26]
  reg  age2_30; // @[DCache.scala 56:26]
  reg  age2_31; // @[DCache.scala 56:26]
  reg [52:0] tag2_0; // @[DCache.scala 57:26]
  reg [52:0] tag2_1; // @[DCache.scala 57:26]
  reg [52:0] tag2_2; // @[DCache.scala 57:26]
  reg [52:0] tag2_3; // @[DCache.scala 57:26]
  reg [52:0] tag2_4; // @[DCache.scala 57:26]
  reg [52:0] tag2_5; // @[DCache.scala 57:26]
  reg [52:0] tag2_6; // @[DCache.scala 57:26]
  reg [52:0] tag2_7; // @[DCache.scala 57:26]
  reg [52:0] tag2_8; // @[DCache.scala 57:26]
  reg [52:0] tag2_9; // @[DCache.scala 57:26]
  reg [52:0] tag2_10; // @[DCache.scala 57:26]
  reg [52:0] tag2_11; // @[DCache.scala 57:26]
  reg [52:0] tag2_12; // @[DCache.scala 57:26]
  reg [52:0] tag2_13; // @[DCache.scala 57:26]
  reg [52:0] tag2_14; // @[DCache.scala 57:26]
  reg [52:0] tag2_15; // @[DCache.scala 57:26]
  reg [52:0] tag2_16; // @[DCache.scala 57:26]
  reg [52:0] tag2_17; // @[DCache.scala 57:26]
  reg [52:0] tag2_18; // @[DCache.scala 57:26]
  reg [52:0] tag2_19; // @[DCache.scala 57:26]
  reg [52:0] tag2_20; // @[DCache.scala 57:26]
  reg [52:0] tag2_21; // @[DCache.scala 57:26]
  reg [52:0] tag2_22; // @[DCache.scala 57:26]
  reg [52:0] tag2_23; // @[DCache.scala 57:26]
  reg [52:0] tag2_24; // @[DCache.scala 57:26]
  reg [52:0] tag2_25; // @[DCache.scala 57:26]
  reg [52:0] tag2_26; // @[DCache.scala 57:26]
  reg [52:0] tag2_27; // @[DCache.scala 57:26]
  reg [52:0] tag2_28; // @[DCache.scala 57:26]
  reg [52:0] tag2_29; // @[DCache.scala 57:26]
  reg [52:0] tag2_30; // @[DCache.scala 57:26]
  reg [52:0] tag2_31; // @[DCache.scala 57:26]
  reg [511:0] block2_0; // @[DCache.scala 58:26]
  reg [511:0] block2_1; // @[DCache.scala 58:26]
  reg [511:0] block2_2; // @[DCache.scala 58:26]
  reg [511:0] block2_3; // @[DCache.scala 58:26]
  reg [511:0] block2_4; // @[DCache.scala 58:26]
  reg [511:0] block2_5; // @[DCache.scala 58:26]
  reg [511:0] block2_6; // @[DCache.scala 58:26]
  reg [511:0] block2_7; // @[DCache.scala 58:26]
  reg [511:0] block2_8; // @[DCache.scala 58:26]
  reg [511:0] block2_9; // @[DCache.scala 58:26]
  reg [511:0] block2_10; // @[DCache.scala 58:26]
  reg [511:0] block2_11; // @[DCache.scala 58:26]
  reg [511:0] block2_12; // @[DCache.scala 58:26]
  reg [511:0] block2_13; // @[DCache.scala 58:26]
  reg [511:0] block2_14; // @[DCache.scala 58:26]
  reg [511:0] block2_15; // @[DCache.scala 58:26]
  reg [511:0] block2_16; // @[DCache.scala 58:26]
  reg [511:0] block2_17; // @[DCache.scala 58:26]
  reg [511:0] block2_18; // @[DCache.scala 58:26]
  reg [511:0] block2_19; // @[DCache.scala 58:26]
  reg [511:0] block2_20; // @[DCache.scala 58:26]
  reg [511:0] block2_21; // @[DCache.scala 58:26]
  reg [511:0] block2_22; // @[DCache.scala 58:26]
  reg [511:0] block2_23; // @[DCache.scala 58:26]
  reg [511:0] block2_24; // @[DCache.scala 58:26]
  reg [511:0] block2_25; // @[DCache.scala 58:26]
  reg [511:0] block2_26; // @[DCache.scala 58:26]
  reg [511:0] block2_27; // @[DCache.scala 58:26]
  reg [511:0] block2_28; // @[DCache.scala 58:26]
  reg [511:0] block2_29; // @[DCache.scala 58:26]
  reg [511:0] block2_30; // @[DCache.scala 58:26]
  reg [511:0] block2_31; // @[DCache.scala 58:26]
  wire [52:0] _GEN_5 = 5'h1 == index_addr ? tag1_1 : tag1_0; // @[DCache.scala 60:28 DCache.scala 60:28]
  wire [52:0] _GEN_6 = 5'h2 == index_addr ? tag1_2 : _GEN_5; // @[DCache.scala 60:28 DCache.scala 60:28]
  wire [52:0] _GEN_7 = 5'h3 == index_addr ? tag1_3 : _GEN_6; // @[DCache.scala 60:28 DCache.scala 60:28]
  wire [52:0] _GEN_8 = 5'h4 == index_addr ? tag1_4 : _GEN_7; // @[DCache.scala 60:28 DCache.scala 60:28]
  wire [52:0] _GEN_9 = 5'h5 == index_addr ? tag1_5 : _GEN_8; // @[DCache.scala 60:28 DCache.scala 60:28]
  wire [52:0] _GEN_10 = 5'h6 == index_addr ? tag1_6 : _GEN_9; // @[DCache.scala 60:28 DCache.scala 60:28]
  wire [52:0] _GEN_11 = 5'h7 == index_addr ? tag1_7 : _GEN_10; // @[DCache.scala 60:28 DCache.scala 60:28]
  wire [52:0] _GEN_12 = 5'h8 == index_addr ? tag1_8 : _GEN_11; // @[DCache.scala 60:28 DCache.scala 60:28]
  wire [52:0] _GEN_13 = 5'h9 == index_addr ? tag1_9 : _GEN_12; // @[DCache.scala 60:28 DCache.scala 60:28]
  wire [52:0] _GEN_14 = 5'ha == index_addr ? tag1_10 : _GEN_13; // @[DCache.scala 60:28 DCache.scala 60:28]
  wire [52:0] _GEN_15 = 5'hb == index_addr ? tag1_11 : _GEN_14; // @[DCache.scala 60:28 DCache.scala 60:28]
  wire [52:0] _GEN_16 = 5'hc == index_addr ? tag1_12 : _GEN_15; // @[DCache.scala 60:28 DCache.scala 60:28]
  wire [52:0] _GEN_17 = 5'hd == index_addr ? tag1_13 : _GEN_16; // @[DCache.scala 60:28 DCache.scala 60:28]
  wire [52:0] _GEN_18 = 5'he == index_addr ? tag1_14 : _GEN_17; // @[DCache.scala 60:28 DCache.scala 60:28]
  wire [52:0] _GEN_19 = 5'hf == index_addr ? tag1_15 : _GEN_18; // @[DCache.scala 60:28 DCache.scala 60:28]
  wire [52:0] _GEN_20 = 5'h10 == index_addr ? tag1_16 : _GEN_19; // @[DCache.scala 60:28 DCache.scala 60:28]
  wire [52:0] _GEN_21 = 5'h11 == index_addr ? tag1_17 : _GEN_20; // @[DCache.scala 60:28 DCache.scala 60:28]
  wire [52:0] _GEN_22 = 5'h12 == index_addr ? tag1_18 : _GEN_21; // @[DCache.scala 60:28 DCache.scala 60:28]
  wire [52:0] _GEN_23 = 5'h13 == index_addr ? tag1_19 : _GEN_22; // @[DCache.scala 60:28 DCache.scala 60:28]
  wire [52:0] _GEN_24 = 5'h14 == index_addr ? tag1_20 : _GEN_23; // @[DCache.scala 60:28 DCache.scala 60:28]
  wire [52:0] _GEN_25 = 5'h15 == index_addr ? tag1_21 : _GEN_24; // @[DCache.scala 60:28 DCache.scala 60:28]
  wire [52:0] _GEN_26 = 5'h16 == index_addr ? tag1_22 : _GEN_25; // @[DCache.scala 60:28 DCache.scala 60:28]
  wire [52:0] _GEN_27 = 5'h17 == index_addr ? tag1_23 : _GEN_26; // @[DCache.scala 60:28 DCache.scala 60:28]
  wire [52:0] _GEN_28 = 5'h18 == index_addr ? tag1_24 : _GEN_27; // @[DCache.scala 60:28 DCache.scala 60:28]
  wire [52:0] _GEN_29 = 5'h19 == index_addr ? tag1_25 : _GEN_28; // @[DCache.scala 60:28 DCache.scala 60:28]
  wire [52:0] _GEN_30 = 5'h1a == index_addr ? tag1_26 : _GEN_29; // @[DCache.scala 60:28 DCache.scala 60:28]
  wire [52:0] _GEN_31 = 5'h1b == index_addr ? tag1_27 : _GEN_30; // @[DCache.scala 60:28 DCache.scala 60:28]
  wire [52:0] _GEN_32 = 5'h1c == index_addr ? tag1_28 : _GEN_31; // @[DCache.scala 60:28 DCache.scala 60:28]
  wire [52:0] _GEN_33 = 5'h1d == index_addr ? tag1_29 : _GEN_32; // @[DCache.scala 60:28 DCache.scala 60:28]
  wire [52:0] _GEN_34 = 5'h1e == index_addr ? tag1_30 : _GEN_33; // @[DCache.scala 60:28 DCache.scala 60:28]
  wire [52:0] _GEN_35 = 5'h1f == index_addr ? tag1_31 : _GEN_34; // @[DCache.scala 60:28 DCache.scala 60:28]
  wire  _GEN_37 = 5'h1 == index_addr ? v1_1 : v1_0; // @[DCache.scala 60:67 DCache.scala 60:67]
  wire  _GEN_38 = 5'h2 == index_addr ? v1_2 : _GEN_37; // @[DCache.scala 60:67 DCache.scala 60:67]
  wire  _GEN_39 = 5'h3 == index_addr ? v1_3 : _GEN_38; // @[DCache.scala 60:67 DCache.scala 60:67]
  wire  _GEN_40 = 5'h4 == index_addr ? v1_4 : _GEN_39; // @[DCache.scala 60:67 DCache.scala 60:67]
  wire  _GEN_41 = 5'h5 == index_addr ? v1_5 : _GEN_40; // @[DCache.scala 60:67 DCache.scala 60:67]
  wire  _GEN_42 = 5'h6 == index_addr ? v1_6 : _GEN_41; // @[DCache.scala 60:67 DCache.scala 60:67]
  wire  _GEN_43 = 5'h7 == index_addr ? v1_7 : _GEN_42; // @[DCache.scala 60:67 DCache.scala 60:67]
  wire  _GEN_44 = 5'h8 == index_addr ? v1_8 : _GEN_43; // @[DCache.scala 60:67 DCache.scala 60:67]
  wire  _GEN_45 = 5'h9 == index_addr ? v1_9 : _GEN_44; // @[DCache.scala 60:67 DCache.scala 60:67]
  wire  _GEN_46 = 5'ha == index_addr ? v1_10 : _GEN_45; // @[DCache.scala 60:67 DCache.scala 60:67]
  wire  _GEN_47 = 5'hb == index_addr ? v1_11 : _GEN_46; // @[DCache.scala 60:67 DCache.scala 60:67]
  wire  _GEN_48 = 5'hc == index_addr ? v1_12 : _GEN_47; // @[DCache.scala 60:67 DCache.scala 60:67]
  wire  _GEN_49 = 5'hd == index_addr ? v1_13 : _GEN_48; // @[DCache.scala 60:67 DCache.scala 60:67]
  wire  _GEN_50 = 5'he == index_addr ? v1_14 : _GEN_49; // @[DCache.scala 60:67 DCache.scala 60:67]
  wire  _GEN_51 = 5'hf == index_addr ? v1_15 : _GEN_50; // @[DCache.scala 60:67 DCache.scala 60:67]
  wire  _GEN_52 = 5'h10 == index_addr ? v1_16 : _GEN_51; // @[DCache.scala 60:67 DCache.scala 60:67]
  wire  _GEN_53 = 5'h11 == index_addr ? v1_17 : _GEN_52; // @[DCache.scala 60:67 DCache.scala 60:67]
  wire  _GEN_54 = 5'h12 == index_addr ? v1_18 : _GEN_53; // @[DCache.scala 60:67 DCache.scala 60:67]
  wire  _GEN_55 = 5'h13 == index_addr ? v1_19 : _GEN_54; // @[DCache.scala 60:67 DCache.scala 60:67]
  wire  _GEN_56 = 5'h14 == index_addr ? v1_20 : _GEN_55; // @[DCache.scala 60:67 DCache.scala 60:67]
  wire  _GEN_57 = 5'h15 == index_addr ? v1_21 : _GEN_56; // @[DCache.scala 60:67 DCache.scala 60:67]
  wire  _GEN_58 = 5'h16 == index_addr ? v1_22 : _GEN_57; // @[DCache.scala 60:67 DCache.scala 60:67]
  wire  _GEN_59 = 5'h17 == index_addr ? v1_23 : _GEN_58; // @[DCache.scala 60:67 DCache.scala 60:67]
  wire  _GEN_60 = 5'h18 == index_addr ? v1_24 : _GEN_59; // @[DCache.scala 60:67 DCache.scala 60:67]
  wire  _GEN_61 = 5'h19 == index_addr ? v1_25 : _GEN_60; // @[DCache.scala 60:67 DCache.scala 60:67]
  wire  _GEN_62 = 5'h1a == index_addr ? v1_26 : _GEN_61; // @[DCache.scala 60:67 DCache.scala 60:67]
  wire  _GEN_63 = 5'h1b == index_addr ? v1_27 : _GEN_62; // @[DCache.scala 60:67 DCache.scala 60:67]
  wire  _GEN_64 = 5'h1c == index_addr ? v1_28 : _GEN_63; // @[DCache.scala 60:67 DCache.scala 60:67]
  wire  _GEN_65 = 5'h1d == index_addr ? v1_29 : _GEN_64; // @[DCache.scala 60:67 DCache.scala 60:67]
  wire  _GEN_66 = 5'h1e == index_addr ? v1_30 : _GEN_65; // @[DCache.scala 60:67 DCache.scala 60:67]
  wire  _GEN_67 = 5'h1f == index_addr ? v1_31 : _GEN_66; // @[DCache.scala 60:67 DCache.scala 60:67]
  wire  hit1 = tag_addr == _GEN_35 & _GEN_67; // @[DCache.scala 60:49]
  wire [52:0] _GEN_69 = 5'h1 == index_addr ? tag2_1 : tag2_0; // @[DCache.scala 61:28 DCache.scala 61:28]
  wire [52:0] _GEN_70 = 5'h2 == index_addr ? tag2_2 : _GEN_69; // @[DCache.scala 61:28 DCache.scala 61:28]
  wire [52:0] _GEN_71 = 5'h3 == index_addr ? tag2_3 : _GEN_70; // @[DCache.scala 61:28 DCache.scala 61:28]
  wire [52:0] _GEN_72 = 5'h4 == index_addr ? tag2_4 : _GEN_71; // @[DCache.scala 61:28 DCache.scala 61:28]
  wire [52:0] _GEN_73 = 5'h5 == index_addr ? tag2_5 : _GEN_72; // @[DCache.scala 61:28 DCache.scala 61:28]
  wire [52:0] _GEN_74 = 5'h6 == index_addr ? tag2_6 : _GEN_73; // @[DCache.scala 61:28 DCache.scala 61:28]
  wire [52:0] _GEN_75 = 5'h7 == index_addr ? tag2_7 : _GEN_74; // @[DCache.scala 61:28 DCache.scala 61:28]
  wire [52:0] _GEN_76 = 5'h8 == index_addr ? tag2_8 : _GEN_75; // @[DCache.scala 61:28 DCache.scala 61:28]
  wire [52:0] _GEN_77 = 5'h9 == index_addr ? tag2_9 : _GEN_76; // @[DCache.scala 61:28 DCache.scala 61:28]
  wire [52:0] _GEN_78 = 5'ha == index_addr ? tag2_10 : _GEN_77; // @[DCache.scala 61:28 DCache.scala 61:28]
  wire [52:0] _GEN_79 = 5'hb == index_addr ? tag2_11 : _GEN_78; // @[DCache.scala 61:28 DCache.scala 61:28]
  wire [52:0] _GEN_80 = 5'hc == index_addr ? tag2_12 : _GEN_79; // @[DCache.scala 61:28 DCache.scala 61:28]
  wire [52:0] _GEN_81 = 5'hd == index_addr ? tag2_13 : _GEN_80; // @[DCache.scala 61:28 DCache.scala 61:28]
  wire [52:0] _GEN_82 = 5'he == index_addr ? tag2_14 : _GEN_81; // @[DCache.scala 61:28 DCache.scala 61:28]
  wire [52:0] _GEN_83 = 5'hf == index_addr ? tag2_15 : _GEN_82; // @[DCache.scala 61:28 DCache.scala 61:28]
  wire [52:0] _GEN_84 = 5'h10 == index_addr ? tag2_16 : _GEN_83; // @[DCache.scala 61:28 DCache.scala 61:28]
  wire [52:0] _GEN_85 = 5'h11 == index_addr ? tag2_17 : _GEN_84; // @[DCache.scala 61:28 DCache.scala 61:28]
  wire [52:0] _GEN_86 = 5'h12 == index_addr ? tag2_18 : _GEN_85; // @[DCache.scala 61:28 DCache.scala 61:28]
  wire [52:0] _GEN_87 = 5'h13 == index_addr ? tag2_19 : _GEN_86; // @[DCache.scala 61:28 DCache.scala 61:28]
  wire [52:0] _GEN_88 = 5'h14 == index_addr ? tag2_20 : _GEN_87; // @[DCache.scala 61:28 DCache.scala 61:28]
  wire [52:0] _GEN_89 = 5'h15 == index_addr ? tag2_21 : _GEN_88; // @[DCache.scala 61:28 DCache.scala 61:28]
  wire [52:0] _GEN_90 = 5'h16 == index_addr ? tag2_22 : _GEN_89; // @[DCache.scala 61:28 DCache.scala 61:28]
  wire [52:0] _GEN_91 = 5'h17 == index_addr ? tag2_23 : _GEN_90; // @[DCache.scala 61:28 DCache.scala 61:28]
  wire [52:0] _GEN_92 = 5'h18 == index_addr ? tag2_24 : _GEN_91; // @[DCache.scala 61:28 DCache.scala 61:28]
  wire [52:0] _GEN_93 = 5'h19 == index_addr ? tag2_25 : _GEN_92; // @[DCache.scala 61:28 DCache.scala 61:28]
  wire [52:0] _GEN_94 = 5'h1a == index_addr ? tag2_26 : _GEN_93; // @[DCache.scala 61:28 DCache.scala 61:28]
  wire [52:0] _GEN_95 = 5'h1b == index_addr ? tag2_27 : _GEN_94; // @[DCache.scala 61:28 DCache.scala 61:28]
  wire [52:0] _GEN_96 = 5'h1c == index_addr ? tag2_28 : _GEN_95; // @[DCache.scala 61:28 DCache.scala 61:28]
  wire [52:0] _GEN_97 = 5'h1d == index_addr ? tag2_29 : _GEN_96; // @[DCache.scala 61:28 DCache.scala 61:28]
  wire [52:0] _GEN_98 = 5'h1e == index_addr ? tag2_30 : _GEN_97; // @[DCache.scala 61:28 DCache.scala 61:28]
  wire [52:0] _GEN_99 = 5'h1f == index_addr ? tag2_31 : _GEN_98; // @[DCache.scala 61:28 DCache.scala 61:28]
  wire  _GEN_101 = 5'h1 == index_addr ? v2_1 : v2_0; // @[DCache.scala 61:67 DCache.scala 61:67]
  wire  _GEN_102 = 5'h2 == index_addr ? v2_2 : _GEN_101; // @[DCache.scala 61:67 DCache.scala 61:67]
  wire  _GEN_103 = 5'h3 == index_addr ? v2_3 : _GEN_102; // @[DCache.scala 61:67 DCache.scala 61:67]
  wire  _GEN_104 = 5'h4 == index_addr ? v2_4 : _GEN_103; // @[DCache.scala 61:67 DCache.scala 61:67]
  wire  _GEN_105 = 5'h5 == index_addr ? v2_5 : _GEN_104; // @[DCache.scala 61:67 DCache.scala 61:67]
  wire  _GEN_106 = 5'h6 == index_addr ? v2_6 : _GEN_105; // @[DCache.scala 61:67 DCache.scala 61:67]
  wire  _GEN_107 = 5'h7 == index_addr ? v2_7 : _GEN_106; // @[DCache.scala 61:67 DCache.scala 61:67]
  wire  _GEN_108 = 5'h8 == index_addr ? v2_8 : _GEN_107; // @[DCache.scala 61:67 DCache.scala 61:67]
  wire  _GEN_109 = 5'h9 == index_addr ? v2_9 : _GEN_108; // @[DCache.scala 61:67 DCache.scala 61:67]
  wire  _GEN_110 = 5'ha == index_addr ? v2_10 : _GEN_109; // @[DCache.scala 61:67 DCache.scala 61:67]
  wire  _GEN_111 = 5'hb == index_addr ? v2_11 : _GEN_110; // @[DCache.scala 61:67 DCache.scala 61:67]
  wire  _GEN_112 = 5'hc == index_addr ? v2_12 : _GEN_111; // @[DCache.scala 61:67 DCache.scala 61:67]
  wire  _GEN_113 = 5'hd == index_addr ? v2_13 : _GEN_112; // @[DCache.scala 61:67 DCache.scala 61:67]
  wire  _GEN_114 = 5'he == index_addr ? v2_14 : _GEN_113; // @[DCache.scala 61:67 DCache.scala 61:67]
  wire  _GEN_115 = 5'hf == index_addr ? v2_15 : _GEN_114; // @[DCache.scala 61:67 DCache.scala 61:67]
  wire  _GEN_116 = 5'h10 == index_addr ? v2_16 : _GEN_115; // @[DCache.scala 61:67 DCache.scala 61:67]
  wire  _GEN_117 = 5'h11 == index_addr ? v2_17 : _GEN_116; // @[DCache.scala 61:67 DCache.scala 61:67]
  wire  _GEN_118 = 5'h12 == index_addr ? v2_18 : _GEN_117; // @[DCache.scala 61:67 DCache.scala 61:67]
  wire  _GEN_119 = 5'h13 == index_addr ? v2_19 : _GEN_118; // @[DCache.scala 61:67 DCache.scala 61:67]
  wire  _GEN_120 = 5'h14 == index_addr ? v2_20 : _GEN_119; // @[DCache.scala 61:67 DCache.scala 61:67]
  wire  _GEN_121 = 5'h15 == index_addr ? v2_21 : _GEN_120; // @[DCache.scala 61:67 DCache.scala 61:67]
  wire  _GEN_122 = 5'h16 == index_addr ? v2_22 : _GEN_121; // @[DCache.scala 61:67 DCache.scala 61:67]
  wire  _GEN_123 = 5'h17 == index_addr ? v2_23 : _GEN_122; // @[DCache.scala 61:67 DCache.scala 61:67]
  wire  _GEN_124 = 5'h18 == index_addr ? v2_24 : _GEN_123; // @[DCache.scala 61:67 DCache.scala 61:67]
  wire  _GEN_125 = 5'h19 == index_addr ? v2_25 : _GEN_124; // @[DCache.scala 61:67 DCache.scala 61:67]
  wire  _GEN_126 = 5'h1a == index_addr ? v2_26 : _GEN_125; // @[DCache.scala 61:67 DCache.scala 61:67]
  wire  _GEN_127 = 5'h1b == index_addr ? v2_27 : _GEN_126; // @[DCache.scala 61:67 DCache.scala 61:67]
  wire  _GEN_128 = 5'h1c == index_addr ? v2_28 : _GEN_127; // @[DCache.scala 61:67 DCache.scala 61:67]
  wire  _GEN_129 = 5'h1d == index_addr ? v2_29 : _GEN_128; // @[DCache.scala 61:67 DCache.scala 61:67]
  wire  _GEN_130 = 5'h1e == index_addr ? v2_30 : _GEN_129; // @[DCache.scala 61:67 DCache.scala 61:67]
  wire  _GEN_131 = 5'h1f == index_addr ? v2_31 : _GEN_130; // @[DCache.scala 61:67 DCache.scala 61:67]
  wire  hit2 = tag_addr == _GEN_99 & _GEN_131; // @[DCache.scala 61:49]
  wire [8:0] _rdata1_T = {offset_addr, 3'h0}; // @[DCache.scala 62:55]
  wire [511:0] _GEN_133 = 5'h1 == index_addr ? block1_1 : block1_0; // @[DCache.scala 62:39 DCache.scala 62:39]
  wire [511:0] _GEN_134 = 5'h2 == index_addr ? block1_2 : _GEN_133; // @[DCache.scala 62:39 DCache.scala 62:39]
  wire [511:0] _GEN_135 = 5'h3 == index_addr ? block1_3 : _GEN_134; // @[DCache.scala 62:39 DCache.scala 62:39]
  wire [511:0] _GEN_136 = 5'h4 == index_addr ? block1_4 : _GEN_135; // @[DCache.scala 62:39 DCache.scala 62:39]
  wire [511:0] _GEN_137 = 5'h5 == index_addr ? block1_5 : _GEN_136; // @[DCache.scala 62:39 DCache.scala 62:39]
  wire [511:0] _GEN_138 = 5'h6 == index_addr ? block1_6 : _GEN_137; // @[DCache.scala 62:39 DCache.scala 62:39]
  wire [511:0] _GEN_139 = 5'h7 == index_addr ? block1_7 : _GEN_138; // @[DCache.scala 62:39 DCache.scala 62:39]
  wire [511:0] _GEN_140 = 5'h8 == index_addr ? block1_8 : _GEN_139; // @[DCache.scala 62:39 DCache.scala 62:39]
  wire [511:0] _GEN_141 = 5'h9 == index_addr ? block1_9 : _GEN_140; // @[DCache.scala 62:39 DCache.scala 62:39]
  wire [511:0] _GEN_142 = 5'ha == index_addr ? block1_10 : _GEN_141; // @[DCache.scala 62:39 DCache.scala 62:39]
  wire [511:0] _GEN_143 = 5'hb == index_addr ? block1_11 : _GEN_142; // @[DCache.scala 62:39 DCache.scala 62:39]
  wire [511:0] _GEN_144 = 5'hc == index_addr ? block1_12 : _GEN_143; // @[DCache.scala 62:39 DCache.scala 62:39]
  wire [511:0] _GEN_145 = 5'hd == index_addr ? block1_13 : _GEN_144; // @[DCache.scala 62:39 DCache.scala 62:39]
  wire [511:0] _GEN_146 = 5'he == index_addr ? block1_14 : _GEN_145; // @[DCache.scala 62:39 DCache.scala 62:39]
  wire [511:0] _GEN_147 = 5'hf == index_addr ? block1_15 : _GEN_146; // @[DCache.scala 62:39 DCache.scala 62:39]
  wire [511:0] _GEN_148 = 5'h10 == index_addr ? block1_16 : _GEN_147; // @[DCache.scala 62:39 DCache.scala 62:39]
  wire [511:0] _GEN_149 = 5'h11 == index_addr ? block1_17 : _GEN_148; // @[DCache.scala 62:39 DCache.scala 62:39]
  wire [511:0] _GEN_150 = 5'h12 == index_addr ? block1_18 : _GEN_149; // @[DCache.scala 62:39 DCache.scala 62:39]
  wire [511:0] _GEN_151 = 5'h13 == index_addr ? block1_19 : _GEN_150; // @[DCache.scala 62:39 DCache.scala 62:39]
  wire [511:0] _GEN_152 = 5'h14 == index_addr ? block1_20 : _GEN_151; // @[DCache.scala 62:39 DCache.scala 62:39]
  wire [511:0] _GEN_153 = 5'h15 == index_addr ? block1_21 : _GEN_152; // @[DCache.scala 62:39 DCache.scala 62:39]
  wire [511:0] _GEN_154 = 5'h16 == index_addr ? block1_22 : _GEN_153; // @[DCache.scala 62:39 DCache.scala 62:39]
  wire [511:0] _GEN_155 = 5'h17 == index_addr ? block1_23 : _GEN_154; // @[DCache.scala 62:39 DCache.scala 62:39]
  wire [511:0] _GEN_156 = 5'h18 == index_addr ? block1_24 : _GEN_155; // @[DCache.scala 62:39 DCache.scala 62:39]
  wire [511:0] _GEN_157 = 5'h19 == index_addr ? block1_25 : _GEN_156; // @[DCache.scala 62:39 DCache.scala 62:39]
  wire [511:0] _GEN_158 = 5'h1a == index_addr ? block1_26 : _GEN_157; // @[DCache.scala 62:39 DCache.scala 62:39]
  wire [511:0] _GEN_159 = 5'h1b == index_addr ? block1_27 : _GEN_158; // @[DCache.scala 62:39 DCache.scala 62:39]
  wire [511:0] _GEN_160 = 5'h1c == index_addr ? block1_28 : _GEN_159; // @[DCache.scala 62:39 DCache.scala 62:39]
  wire [511:0] _GEN_161 = 5'h1d == index_addr ? block1_29 : _GEN_160; // @[DCache.scala 62:39 DCache.scala 62:39]
  wire [511:0] _GEN_162 = 5'h1e == index_addr ? block1_30 : _GEN_161; // @[DCache.scala 62:39 DCache.scala 62:39]
  wire [511:0] _GEN_163 = 5'h1f == index_addr ? block1_31 : _GEN_162; // @[DCache.scala 62:39 DCache.scala 62:39]
  wire [511:0] _rdata1_T_1 = _GEN_163 >> _rdata1_T; // @[DCache.scala 62:39]
  wire [63:0] rdata1 = _rdata1_T_1[63:0]; // @[DCache.scala 62:61]
  wire [511:0] _GEN_165 = 5'h1 == index_addr ? block2_1 : block2_0; // @[DCache.scala 63:39 DCache.scala 63:39]
  wire [511:0] _GEN_166 = 5'h2 == index_addr ? block2_2 : _GEN_165; // @[DCache.scala 63:39 DCache.scala 63:39]
  wire [511:0] _GEN_167 = 5'h3 == index_addr ? block2_3 : _GEN_166; // @[DCache.scala 63:39 DCache.scala 63:39]
  wire [511:0] _GEN_168 = 5'h4 == index_addr ? block2_4 : _GEN_167; // @[DCache.scala 63:39 DCache.scala 63:39]
  wire [511:0] _GEN_169 = 5'h5 == index_addr ? block2_5 : _GEN_168; // @[DCache.scala 63:39 DCache.scala 63:39]
  wire [511:0] _GEN_170 = 5'h6 == index_addr ? block2_6 : _GEN_169; // @[DCache.scala 63:39 DCache.scala 63:39]
  wire [511:0] _GEN_171 = 5'h7 == index_addr ? block2_7 : _GEN_170; // @[DCache.scala 63:39 DCache.scala 63:39]
  wire [511:0] _GEN_172 = 5'h8 == index_addr ? block2_8 : _GEN_171; // @[DCache.scala 63:39 DCache.scala 63:39]
  wire [511:0] _GEN_173 = 5'h9 == index_addr ? block2_9 : _GEN_172; // @[DCache.scala 63:39 DCache.scala 63:39]
  wire [511:0] _GEN_174 = 5'ha == index_addr ? block2_10 : _GEN_173; // @[DCache.scala 63:39 DCache.scala 63:39]
  wire [511:0] _GEN_175 = 5'hb == index_addr ? block2_11 : _GEN_174; // @[DCache.scala 63:39 DCache.scala 63:39]
  wire [511:0] _GEN_176 = 5'hc == index_addr ? block2_12 : _GEN_175; // @[DCache.scala 63:39 DCache.scala 63:39]
  wire [511:0] _GEN_177 = 5'hd == index_addr ? block2_13 : _GEN_176; // @[DCache.scala 63:39 DCache.scala 63:39]
  wire [511:0] _GEN_178 = 5'he == index_addr ? block2_14 : _GEN_177; // @[DCache.scala 63:39 DCache.scala 63:39]
  wire [511:0] _GEN_179 = 5'hf == index_addr ? block2_15 : _GEN_178; // @[DCache.scala 63:39 DCache.scala 63:39]
  wire [511:0] _GEN_180 = 5'h10 == index_addr ? block2_16 : _GEN_179; // @[DCache.scala 63:39 DCache.scala 63:39]
  wire [511:0] _GEN_181 = 5'h11 == index_addr ? block2_17 : _GEN_180; // @[DCache.scala 63:39 DCache.scala 63:39]
  wire [511:0] _GEN_182 = 5'h12 == index_addr ? block2_18 : _GEN_181; // @[DCache.scala 63:39 DCache.scala 63:39]
  wire [511:0] _GEN_183 = 5'h13 == index_addr ? block2_19 : _GEN_182; // @[DCache.scala 63:39 DCache.scala 63:39]
  wire [511:0] _GEN_184 = 5'h14 == index_addr ? block2_20 : _GEN_183; // @[DCache.scala 63:39 DCache.scala 63:39]
  wire [511:0] _GEN_185 = 5'h15 == index_addr ? block2_21 : _GEN_184; // @[DCache.scala 63:39 DCache.scala 63:39]
  wire [511:0] _GEN_186 = 5'h16 == index_addr ? block2_22 : _GEN_185; // @[DCache.scala 63:39 DCache.scala 63:39]
  wire [511:0] _GEN_187 = 5'h17 == index_addr ? block2_23 : _GEN_186; // @[DCache.scala 63:39 DCache.scala 63:39]
  wire [511:0] _GEN_188 = 5'h18 == index_addr ? block2_24 : _GEN_187; // @[DCache.scala 63:39 DCache.scala 63:39]
  wire [511:0] _GEN_189 = 5'h19 == index_addr ? block2_25 : _GEN_188; // @[DCache.scala 63:39 DCache.scala 63:39]
  wire [511:0] _GEN_190 = 5'h1a == index_addr ? block2_26 : _GEN_189; // @[DCache.scala 63:39 DCache.scala 63:39]
  wire [511:0] _GEN_191 = 5'h1b == index_addr ? block2_27 : _GEN_190; // @[DCache.scala 63:39 DCache.scala 63:39]
  wire [511:0] _GEN_192 = 5'h1c == index_addr ? block2_28 : _GEN_191; // @[DCache.scala 63:39 DCache.scala 63:39]
  wire [511:0] _GEN_193 = 5'h1d == index_addr ? block2_29 : _GEN_192; // @[DCache.scala 63:39 DCache.scala 63:39]
  wire [511:0] _GEN_194 = 5'h1e == index_addr ? block2_30 : _GEN_193; // @[DCache.scala 63:39 DCache.scala 63:39]
  wire [511:0] _GEN_195 = 5'h1f == index_addr ? block2_31 : _GEN_194; // @[DCache.scala 63:39 DCache.scala 63:39]
  wire [511:0] _rdata2_T_1 = _GEN_195 >> _rdata1_T; // @[DCache.scala 63:39]
  wire [63:0] rdata2 = _rdata2_T_1[63:0]; // @[DCache.scala 63:61]
  reg [1:0] state; // @[DCache.scala 66:24]
  wire  hit = hit1 | hit2; // @[DCache.scala 68:28]
  wire [63:0] _rdata_T = hit1 ? rdata1 : 64'h0; // @[DCache.scala 69:44]
  reg  not_en_yet; // @[DCache.scala 71:30]
  wire  _not_en_yet_T = io_dmem_en ? 1'h0 : not_en_yet; // @[DCache.scala 72:27]
  wire  _age1_T = hit1 ^ hit2; // @[DCache.scala 78:35]
  wire  _GEN_197 = 5'h1 == index_addr ? age1_1 : age1_0; // @[DCache.scala 78:28 DCache.scala 78:28]
  wire  _GEN_198 = 5'h2 == index_addr ? age1_2 : _GEN_197; // @[DCache.scala 78:28 DCache.scala 78:28]
  wire  _GEN_199 = 5'h3 == index_addr ? age1_3 : _GEN_198; // @[DCache.scala 78:28 DCache.scala 78:28]
  wire  _GEN_200 = 5'h4 == index_addr ? age1_4 : _GEN_199; // @[DCache.scala 78:28 DCache.scala 78:28]
  wire  _GEN_201 = 5'h5 == index_addr ? age1_5 : _GEN_200; // @[DCache.scala 78:28 DCache.scala 78:28]
  wire  _GEN_202 = 5'h6 == index_addr ? age1_6 : _GEN_201; // @[DCache.scala 78:28 DCache.scala 78:28]
  wire  _GEN_203 = 5'h7 == index_addr ? age1_7 : _GEN_202; // @[DCache.scala 78:28 DCache.scala 78:28]
  wire  _GEN_204 = 5'h8 == index_addr ? age1_8 : _GEN_203; // @[DCache.scala 78:28 DCache.scala 78:28]
  wire  _GEN_205 = 5'h9 == index_addr ? age1_9 : _GEN_204; // @[DCache.scala 78:28 DCache.scala 78:28]
  wire  _GEN_206 = 5'ha == index_addr ? age1_10 : _GEN_205; // @[DCache.scala 78:28 DCache.scala 78:28]
  wire  _GEN_207 = 5'hb == index_addr ? age1_11 : _GEN_206; // @[DCache.scala 78:28 DCache.scala 78:28]
  wire  _GEN_208 = 5'hc == index_addr ? age1_12 : _GEN_207; // @[DCache.scala 78:28 DCache.scala 78:28]
  wire  _GEN_209 = 5'hd == index_addr ? age1_13 : _GEN_208; // @[DCache.scala 78:28 DCache.scala 78:28]
  wire  _GEN_210 = 5'he == index_addr ? age1_14 : _GEN_209; // @[DCache.scala 78:28 DCache.scala 78:28]
  wire  _GEN_211 = 5'hf == index_addr ? age1_15 : _GEN_210; // @[DCache.scala 78:28 DCache.scala 78:28]
  wire  _GEN_212 = 5'h10 == index_addr ? age1_16 : _GEN_211; // @[DCache.scala 78:28 DCache.scala 78:28]
  wire  _GEN_213 = 5'h11 == index_addr ? age1_17 : _GEN_212; // @[DCache.scala 78:28 DCache.scala 78:28]
  wire  _GEN_214 = 5'h12 == index_addr ? age1_18 : _GEN_213; // @[DCache.scala 78:28 DCache.scala 78:28]
  wire  _GEN_215 = 5'h13 == index_addr ? age1_19 : _GEN_214; // @[DCache.scala 78:28 DCache.scala 78:28]
  wire  _GEN_216 = 5'h14 == index_addr ? age1_20 : _GEN_215; // @[DCache.scala 78:28 DCache.scala 78:28]
  wire  _GEN_217 = 5'h15 == index_addr ? age1_21 : _GEN_216; // @[DCache.scala 78:28 DCache.scala 78:28]
  wire  _GEN_218 = 5'h16 == index_addr ? age1_22 : _GEN_217; // @[DCache.scala 78:28 DCache.scala 78:28]
  wire  _GEN_219 = 5'h17 == index_addr ? age1_23 : _GEN_218; // @[DCache.scala 78:28 DCache.scala 78:28]
  wire  _GEN_220 = 5'h18 == index_addr ? age1_24 : _GEN_219; // @[DCache.scala 78:28 DCache.scala 78:28]
  wire  _GEN_221 = 5'h19 == index_addr ? age1_25 : _GEN_220; // @[DCache.scala 78:28 DCache.scala 78:28]
  wire  _GEN_222 = 5'h1a == index_addr ? age1_26 : _GEN_221; // @[DCache.scala 78:28 DCache.scala 78:28]
  wire  _GEN_223 = 5'h1b == index_addr ? age1_27 : _GEN_222; // @[DCache.scala 78:28 DCache.scala 78:28]
  wire  _GEN_224 = 5'h1c == index_addr ? age1_28 : _GEN_223; // @[DCache.scala 78:28 DCache.scala 78:28]
  wire  _GEN_225 = 5'h1d == index_addr ? age1_29 : _GEN_224; // @[DCache.scala 78:28 DCache.scala 78:28]
  wire  _GEN_226 = 5'h1e == index_addr ? age1_30 : _GEN_225; // @[DCache.scala 78:28 DCache.scala 78:28]
  wire  _GEN_227 = 5'h1f == index_addr ? age1_31 : _GEN_226; // @[DCache.scala 78:28 DCache.scala 78:28]
  wire  _GEN_261 = 5'h1 == index_addr ? age2_1 : age2_0; // @[DCache.scala 79:28 DCache.scala 79:28]
  wire  _GEN_262 = 5'h2 == index_addr ? age2_2 : _GEN_261; // @[DCache.scala 79:28 DCache.scala 79:28]
  wire  _GEN_263 = 5'h3 == index_addr ? age2_3 : _GEN_262; // @[DCache.scala 79:28 DCache.scala 79:28]
  wire  _GEN_264 = 5'h4 == index_addr ? age2_4 : _GEN_263; // @[DCache.scala 79:28 DCache.scala 79:28]
  wire  _GEN_265 = 5'h5 == index_addr ? age2_5 : _GEN_264; // @[DCache.scala 79:28 DCache.scala 79:28]
  wire  _GEN_266 = 5'h6 == index_addr ? age2_6 : _GEN_265; // @[DCache.scala 79:28 DCache.scala 79:28]
  wire  _GEN_267 = 5'h7 == index_addr ? age2_7 : _GEN_266; // @[DCache.scala 79:28 DCache.scala 79:28]
  wire  _GEN_268 = 5'h8 == index_addr ? age2_8 : _GEN_267; // @[DCache.scala 79:28 DCache.scala 79:28]
  wire  _GEN_269 = 5'h9 == index_addr ? age2_9 : _GEN_268; // @[DCache.scala 79:28 DCache.scala 79:28]
  wire  _GEN_270 = 5'ha == index_addr ? age2_10 : _GEN_269; // @[DCache.scala 79:28 DCache.scala 79:28]
  wire  _GEN_271 = 5'hb == index_addr ? age2_11 : _GEN_270; // @[DCache.scala 79:28 DCache.scala 79:28]
  wire  _GEN_272 = 5'hc == index_addr ? age2_12 : _GEN_271; // @[DCache.scala 79:28 DCache.scala 79:28]
  wire  _GEN_273 = 5'hd == index_addr ? age2_13 : _GEN_272; // @[DCache.scala 79:28 DCache.scala 79:28]
  wire  _GEN_274 = 5'he == index_addr ? age2_14 : _GEN_273; // @[DCache.scala 79:28 DCache.scala 79:28]
  wire  _GEN_275 = 5'hf == index_addr ? age2_15 : _GEN_274; // @[DCache.scala 79:28 DCache.scala 79:28]
  wire  _GEN_276 = 5'h10 == index_addr ? age2_16 : _GEN_275; // @[DCache.scala 79:28 DCache.scala 79:28]
  wire  _GEN_277 = 5'h11 == index_addr ? age2_17 : _GEN_276; // @[DCache.scala 79:28 DCache.scala 79:28]
  wire  _GEN_278 = 5'h12 == index_addr ? age2_18 : _GEN_277; // @[DCache.scala 79:28 DCache.scala 79:28]
  wire  _GEN_279 = 5'h13 == index_addr ? age2_19 : _GEN_278; // @[DCache.scala 79:28 DCache.scala 79:28]
  wire  _GEN_280 = 5'h14 == index_addr ? age2_20 : _GEN_279; // @[DCache.scala 79:28 DCache.scala 79:28]
  wire  _GEN_281 = 5'h15 == index_addr ? age2_21 : _GEN_280; // @[DCache.scala 79:28 DCache.scala 79:28]
  wire  _GEN_282 = 5'h16 == index_addr ? age2_22 : _GEN_281; // @[DCache.scala 79:28 DCache.scala 79:28]
  wire  _GEN_283 = 5'h17 == index_addr ? age2_23 : _GEN_282; // @[DCache.scala 79:28 DCache.scala 79:28]
  wire  _GEN_284 = 5'h18 == index_addr ? age2_24 : _GEN_283; // @[DCache.scala 79:28 DCache.scala 79:28]
  wire  _GEN_285 = 5'h19 == index_addr ? age2_25 : _GEN_284; // @[DCache.scala 79:28 DCache.scala 79:28]
  wire  _GEN_286 = 5'h1a == index_addr ? age2_26 : _GEN_285; // @[DCache.scala 79:28 DCache.scala 79:28]
  wire  _GEN_287 = 5'h1b == index_addr ? age2_27 : _GEN_286; // @[DCache.scala 79:28 DCache.scala 79:28]
  wire  _GEN_288 = 5'h1c == index_addr ? age2_28 : _GEN_287; // @[DCache.scala 79:28 DCache.scala 79:28]
  wire  _GEN_289 = 5'h1d == index_addr ? age2_29 : _GEN_288; // @[DCache.scala 79:28 DCache.scala 79:28]
  wire  _GEN_290 = 5'h1e == index_addr ? age2_30 : _GEN_289; // @[DCache.scala 79:28 DCache.scala 79:28]
  wire  _GEN_291 = 5'h1f == index_addr ? age2_31 : _GEN_290; // @[DCache.scala 79:28 DCache.scala 79:28]
  wire [1:0] age = {_GEN_291,_GEN_227}; // @[Cat.scala 30:58]
  wire  updateway2 = age == 2'h1; // @[DCache.scala 83:27]
  wire  updateway1 = ~updateway2; // @[DCache.scala 84:23]
  wire  miss = ~hit; // @[DCache.scala 85:23]
  wire  _GEN_325 = 5'h1 == index_addr ? d1_1 : d1_0; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_326 = 5'h2 == index_addr ? d1_2 : _GEN_325; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_327 = 5'h3 == index_addr ? d1_3 : _GEN_326; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_328 = 5'h4 == index_addr ? d1_4 : _GEN_327; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_329 = 5'h5 == index_addr ? d1_5 : _GEN_328; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_330 = 5'h6 == index_addr ? d1_6 : _GEN_329; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_331 = 5'h7 == index_addr ? d1_7 : _GEN_330; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_332 = 5'h8 == index_addr ? d1_8 : _GEN_331; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_333 = 5'h9 == index_addr ? d1_9 : _GEN_332; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_334 = 5'ha == index_addr ? d1_10 : _GEN_333; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_335 = 5'hb == index_addr ? d1_11 : _GEN_334; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_336 = 5'hc == index_addr ? d1_12 : _GEN_335; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_337 = 5'hd == index_addr ? d1_13 : _GEN_336; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_338 = 5'he == index_addr ? d1_14 : _GEN_337; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_339 = 5'hf == index_addr ? d1_15 : _GEN_338; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_340 = 5'h10 == index_addr ? d1_16 : _GEN_339; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_341 = 5'h11 == index_addr ? d1_17 : _GEN_340; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_342 = 5'h12 == index_addr ? d1_18 : _GEN_341; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_343 = 5'h13 == index_addr ? d1_19 : _GEN_342; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_344 = 5'h14 == index_addr ? d1_20 : _GEN_343; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_345 = 5'h15 == index_addr ? d1_21 : _GEN_344; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_346 = 5'h16 == index_addr ? d1_22 : _GEN_345; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_347 = 5'h17 == index_addr ? d1_23 : _GEN_346; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_348 = 5'h18 == index_addr ? d1_24 : _GEN_347; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_349 = 5'h19 == index_addr ? d1_25 : _GEN_348; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_350 = 5'h1a == index_addr ? d1_26 : _GEN_349; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_351 = 5'h1b == index_addr ? d1_27 : _GEN_350; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_352 = 5'h1c == index_addr ? d1_28 : _GEN_351; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_353 = 5'h1d == index_addr ? d1_29 : _GEN_352; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_354 = 5'h1e == index_addr ? d1_30 : _GEN_353; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_355 = 5'h1f == index_addr ? d1_31 : _GEN_354; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_357 = 5'h1 == index_addr ? d2_1 : d2_0; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_358 = 5'h2 == index_addr ? d2_2 : _GEN_357; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_359 = 5'h3 == index_addr ? d2_3 : _GEN_358; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_360 = 5'h4 == index_addr ? d2_4 : _GEN_359; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_361 = 5'h5 == index_addr ? d2_5 : _GEN_360; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_362 = 5'h6 == index_addr ? d2_6 : _GEN_361; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_363 = 5'h7 == index_addr ? d2_7 : _GEN_362; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_364 = 5'h8 == index_addr ? d2_8 : _GEN_363; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_365 = 5'h9 == index_addr ? d2_9 : _GEN_364; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_366 = 5'ha == index_addr ? d2_10 : _GEN_365; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_367 = 5'hb == index_addr ? d2_11 : _GEN_366; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_368 = 5'hc == index_addr ? d2_12 : _GEN_367; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_369 = 5'hd == index_addr ? d2_13 : _GEN_368; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_370 = 5'he == index_addr ? d2_14 : _GEN_369; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_371 = 5'hf == index_addr ? d2_15 : _GEN_370; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_372 = 5'h10 == index_addr ? d2_16 : _GEN_371; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_373 = 5'h11 == index_addr ? d2_17 : _GEN_372; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_374 = 5'h12 == index_addr ? d2_18 : _GEN_373; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_375 = 5'h13 == index_addr ? d2_19 : _GEN_374; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_376 = 5'h14 == index_addr ? d2_20 : _GEN_375; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_377 = 5'h15 == index_addr ? d2_21 : _GEN_376; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_378 = 5'h16 == index_addr ? d2_22 : _GEN_377; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_379 = 5'h17 == index_addr ? d2_23 : _GEN_378; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_380 = 5'h18 == index_addr ? d2_24 : _GEN_379; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_381 = 5'h19 == index_addr ? d2_25 : _GEN_380; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_382 = 5'h1a == index_addr ? d2_26 : _GEN_381; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_383 = 5'h1b == index_addr ? d2_27 : _GEN_382; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_384 = 5'h1c == index_addr ? d2_28 : _GEN_383; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_385 = 5'h1d == index_addr ? d2_29 : _GEN_384; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_386 = 5'h1e == index_addr ? d2_30 : _GEN_385; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  _GEN_387 = 5'h1f == index_addr ? d2_31 : _GEN_386; // @[DCache.scala 86:26 DCache.scala 86:26]
  wire  dirty = updateway1 ? _GEN_355 : _GEN_387; // @[DCache.scala 86:26]
  wire  _T = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_3 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_4 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_390 = io_axi_rvalid ? 2'h0 : state; // @[DCache.scala 97:33 DCache.scala 97:40 DCache.scala 66:24]
  wire  update = state == 2'h2 & io_axi_rvalid; // @[DCache.scala 103:39]
  wire  way1write = hit1 & op; // @[DCache.scala 104:26]
  wire  way2write = hit2 & op; // @[DCache.scala 105:26]
  wire  _d1_T = update & updateway1; // @[DCache.scala 106:34]
  wire  _d2_T = update & updateway2; // @[DCache.scala 107:34]
  wire [7:0] mask64_hi_hi_hi_lo = wm[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] mask64_hi_hi_lo = wm[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] mask64_hi_lo_hi = wm[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] mask64_hi_lo_lo = wm[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] mask64_lo_hi_hi = wm[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] mask64_lo_hi_lo = wm[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] mask64_lo_lo_hi = wm[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] mask64_lo_lo_lo = wm[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [511:0] mask64 = {448'h0,mask64_hi_hi_hi_lo,mask64_hi_hi_lo,mask64_hi_lo_hi,mask64_hi_lo_lo,mask64_lo_hi_hi,
    mask64_lo_hi_lo,mask64_lo_lo_hi,mask64_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [8:0] _blockmask_T_1 = {offset_addr[5:3], 6'h0}; // @[DCache.scala 112:52]
  wire [1022:0] _GEN_650 = {{511'd0}, mask64}; // @[DCache.scala 112:29]
  wire [1022:0] _blockmask_T_2 = _GEN_650 << _blockmask_T_1; // @[DCache.scala 112:29]
  wire [511:0] blockmask = _blockmask_T_2[511:0]; // @[DCache.scala 112:58]
  wire [574:0] _GEN_651 = {{511'd0}, wdata}; // @[DCache.scala 113:29]
  wire [574:0] _blockwdata_T_2 = _GEN_651 << _blockmask_T_1; // @[DCache.scala 113:29]
  wire [511:0] blockwdata = _blockwdata_T_2[511:0]; // @[DCache.scala 113:58]
  wire [511:0] _block1_after_write_T = ~blockmask; // @[DCache.scala 114:53]
  wire [511:0] _block1_after_write_T_1 = _GEN_163 & _block1_after_write_T; // @[DCache.scala 114:50]
  wire [511:0] _block1_after_write_T_2 = blockmask & blockwdata; // @[DCache.scala 114:79]
  wire [511:0] block1_after_write = _block1_after_write_T_1 | _block1_after_write_T_2; // @[DCache.scala 114:66]
  wire [511:0] _block2_after_write_T_1 = _GEN_195 & _block1_after_write_T; // @[DCache.scala 115:50]
  wire [511:0] block2_after_write = _block2_after_write_T_1 | _block1_after_write_T_2; // @[DCache.scala 115:66]
  wire [52:0] io_axi_waddr_hi_hi = updateway1 ? _GEN_35 : _GEN_99; // @[DCache.scala 129:31]
  wire [57:0] io_axi_waddr_hi = {io_axi_waddr_hi_hi,index_addr}; // @[Cat.scala 30:58]
  assign io_dmem_ok = (hit | not_en_yet) & state == 2'h0; // @[DCache.scala 75:44]
  assign io_dmem_rdata = hit2 ? rdata2 : _rdata_T; // @[DCache.scala 69:26]
  assign io_axi_req = state == 2'h2; // @[DCache.scala 126:30]
  assign io_axi_raddr = addr & 64'hffffffffffffffc0; // @[DCache.scala 127:29]
  assign io_axi_weq = state == 2'h1; // @[DCache.scala 128:30]
  assign io_axi_waddr = {io_axi_waddr_hi,6'h0}; // @[Cat.scala 30:58]
  assign io_axi_wdata = updateway1 ? _GEN_163 : _GEN_195; // @[DCache.scala 130:27]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 27:20]
      op <= 1'h0; // @[Reg.scala 27:20]
    end else if (_op_T) begin // @[Reg.scala 28:19]
      op <= io_dmem_op; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      addr <= 64'h0; // @[Reg.scala 27:20]
    end else if (_op_T) begin // @[Reg.scala 28:19]
      addr <= io_dmem_addr; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      wdata <= 64'h0; // @[Reg.scala 27:20]
    end else if (_op_T) begin // @[Reg.scala 28:19]
      wdata <= io_dmem_wdata; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      wm <= 8'h0; // @[Reg.scala 27:20]
    end else if (_op_T) begin // @[Reg.scala 28:19]
      wm <= io_dmem_wmask; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[DCache.scala 49:26]
      v1_0 <= 1'h0; // @[DCache.scala 49:26]
    end else if (5'h0 == index_addr) begin // @[DCache.scala 120:26]
      v1_0 <= _d1_T | _GEN_67; // @[DCache.scala 120:26]
    end
    if (reset) begin // @[DCache.scala 49:26]
      v1_1 <= 1'h0; // @[DCache.scala 49:26]
    end else if (5'h1 == index_addr) begin // @[DCache.scala 120:26]
      v1_1 <= _d1_T | _GEN_67; // @[DCache.scala 120:26]
    end
    if (reset) begin // @[DCache.scala 49:26]
      v1_2 <= 1'h0; // @[DCache.scala 49:26]
    end else if (5'h2 == index_addr) begin // @[DCache.scala 120:26]
      v1_2 <= _d1_T | _GEN_67; // @[DCache.scala 120:26]
    end
    if (reset) begin // @[DCache.scala 49:26]
      v1_3 <= 1'h0; // @[DCache.scala 49:26]
    end else if (5'h3 == index_addr) begin // @[DCache.scala 120:26]
      v1_3 <= _d1_T | _GEN_67; // @[DCache.scala 120:26]
    end
    if (reset) begin // @[DCache.scala 49:26]
      v1_4 <= 1'h0; // @[DCache.scala 49:26]
    end else if (5'h4 == index_addr) begin // @[DCache.scala 120:26]
      v1_4 <= _d1_T | _GEN_67; // @[DCache.scala 120:26]
    end
    if (reset) begin // @[DCache.scala 49:26]
      v1_5 <= 1'h0; // @[DCache.scala 49:26]
    end else if (5'h5 == index_addr) begin // @[DCache.scala 120:26]
      v1_5 <= _d1_T | _GEN_67; // @[DCache.scala 120:26]
    end
    if (reset) begin // @[DCache.scala 49:26]
      v1_6 <= 1'h0; // @[DCache.scala 49:26]
    end else if (5'h6 == index_addr) begin // @[DCache.scala 120:26]
      v1_6 <= _d1_T | _GEN_67; // @[DCache.scala 120:26]
    end
    if (reset) begin // @[DCache.scala 49:26]
      v1_7 <= 1'h0; // @[DCache.scala 49:26]
    end else if (5'h7 == index_addr) begin // @[DCache.scala 120:26]
      v1_7 <= _d1_T | _GEN_67; // @[DCache.scala 120:26]
    end
    if (reset) begin // @[DCache.scala 49:26]
      v1_8 <= 1'h0; // @[DCache.scala 49:26]
    end else if (5'h8 == index_addr) begin // @[DCache.scala 120:26]
      v1_8 <= _d1_T | _GEN_67; // @[DCache.scala 120:26]
    end
    if (reset) begin // @[DCache.scala 49:26]
      v1_9 <= 1'h0; // @[DCache.scala 49:26]
    end else if (5'h9 == index_addr) begin // @[DCache.scala 120:26]
      v1_9 <= _d1_T | _GEN_67; // @[DCache.scala 120:26]
    end
    if (reset) begin // @[DCache.scala 49:26]
      v1_10 <= 1'h0; // @[DCache.scala 49:26]
    end else if (5'ha == index_addr) begin // @[DCache.scala 120:26]
      v1_10 <= _d1_T | _GEN_67; // @[DCache.scala 120:26]
    end
    if (reset) begin // @[DCache.scala 49:26]
      v1_11 <= 1'h0; // @[DCache.scala 49:26]
    end else if (5'hb == index_addr) begin // @[DCache.scala 120:26]
      v1_11 <= _d1_T | _GEN_67; // @[DCache.scala 120:26]
    end
    if (reset) begin // @[DCache.scala 49:26]
      v1_12 <= 1'h0; // @[DCache.scala 49:26]
    end else if (5'hc == index_addr) begin // @[DCache.scala 120:26]
      v1_12 <= _d1_T | _GEN_67; // @[DCache.scala 120:26]
    end
    if (reset) begin // @[DCache.scala 49:26]
      v1_13 <= 1'h0; // @[DCache.scala 49:26]
    end else if (5'hd == index_addr) begin // @[DCache.scala 120:26]
      v1_13 <= _d1_T | _GEN_67; // @[DCache.scala 120:26]
    end
    if (reset) begin // @[DCache.scala 49:26]
      v1_14 <= 1'h0; // @[DCache.scala 49:26]
    end else if (5'he == index_addr) begin // @[DCache.scala 120:26]
      v1_14 <= _d1_T | _GEN_67; // @[DCache.scala 120:26]
    end
    if (reset) begin // @[DCache.scala 49:26]
      v1_15 <= 1'h0; // @[DCache.scala 49:26]
    end else if (5'hf == index_addr) begin // @[DCache.scala 120:26]
      v1_15 <= _d1_T | _GEN_67; // @[DCache.scala 120:26]
    end
    if (reset) begin // @[DCache.scala 49:26]
      v1_16 <= 1'h0; // @[DCache.scala 49:26]
    end else if (5'h10 == index_addr) begin // @[DCache.scala 120:26]
      v1_16 <= _d1_T | _GEN_67; // @[DCache.scala 120:26]
    end
    if (reset) begin // @[DCache.scala 49:26]
      v1_17 <= 1'h0; // @[DCache.scala 49:26]
    end else if (5'h11 == index_addr) begin // @[DCache.scala 120:26]
      v1_17 <= _d1_T | _GEN_67; // @[DCache.scala 120:26]
    end
    if (reset) begin // @[DCache.scala 49:26]
      v1_18 <= 1'h0; // @[DCache.scala 49:26]
    end else if (5'h12 == index_addr) begin // @[DCache.scala 120:26]
      v1_18 <= _d1_T | _GEN_67; // @[DCache.scala 120:26]
    end
    if (reset) begin // @[DCache.scala 49:26]
      v1_19 <= 1'h0; // @[DCache.scala 49:26]
    end else if (5'h13 == index_addr) begin // @[DCache.scala 120:26]
      v1_19 <= _d1_T | _GEN_67; // @[DCache.scala 120:26]
    end
    if (reset) begin // @[DCache.scala 49:26]
      v1_20 <= 1'h0; // @[DCache.scala 49:26]
    end else if (5'h14 == index_addr) begin // @[DCache.scala 120:26]
      v1_20 <= _d1_T | _GEN_67; // @[DCache.scala 120:26]
    end
    if (reset) begin // @[DCache.scala 49:26]
      v1_21 <= 1'h0; // @[DCache.scala 49:26]
    end else if (5'h15 == index_addr) begin // @[DCache.scala 120:26]
      v1_21 <= _d1_T | _GEN_67; // @[DCache.scala 120:26]
    end
    if (reset) begin // @[DCache.scala 49:26]
      v1_22 <= 1'h0; // @[DCache.scala 49:26]
    end else if (5'h16 == index_addr) begin // @[DCache.scala 120:26]
      v1_22 <= _d1_T | _GEN_67; // @[DCache.scala 120:26]
    end
    if (reset) begin // @[DCache.scala 49:26]
      v1_23 <= 1'h0; // @[DCache.scala 49:26]
    end else if (5'h17 == index_addr) begin // @[DCache.scala 120:26]
      v1_23 <= _d1_T | _GEN_67; // @[DCache.scala 120:26]
    end
    if (reset) begin // @[DCache.scala 49:26]
      v1_24 <= 1'h0; // @[DCache.scala 49:26]
    end else if (5'h18 == index_addr) begin // @[DCache.scala 120:26]
      v1_24 <= _d1_T | _GEN_67; // @[DCache.scala 120:26]
    end
    if (reset) begin // @[DCache.scala 49:26]
      v1_25 <= 1'h0; // @[DCache.scala 49:26]
    end else if (5'h19 == index_addr) begin // @[DCache.scala 120:26]
      v1_25 <= _d1_T | _GEN_67; // @[DCache.scala 120:26]
    end
    if (reset) begin // @[DCache.scala 49:26]
      v1_26 <= 1'h0; // @[DCache.scala 49:26]
    end else if (5'h1a == index_addr) begin // @[DCache.scala 120:26]
      v1_26 <= _d1_T | _GEN_67; // @[DCache.scala 120:26]
    end
    if (reset) begin // @[DCache.scala 49:26]
      v1_27 <= 1'h0; // @[DCache.scala 49:26]
    end else if (5'h1b == index_addr) begin // @[DCache.scala 120:26]
      v1_27 <= _d1_T | _GEN_67; // @[DCache.scala 120:26]
    end
    if (reset) begin // @[DCache.scala 49:26]
      v1_28 <= 1'h0; // @[DCache.scala 49:26]
    end else if (5'h1c == index_addr) begin // @[DCache.scala 120:26]
      v1_28 <= _d1_T | _GEN_67; // @[DCache.scala 120:26]
    end
    if (reset) begin // @[DCache.scala 49:26]
      v1_29 <= 1'h0; // @[DCache.scala 49:26]
    end else if (5'h1d == index_addr) begin // @[DCache.scala 120:26]
      v1_29 <= _d1_T | _GEN_67; // @[DCache.scala 120:26]
    end
    if (reset) begin // @[DCache.scala 49:26]
      v1_30 <= 1'h0; // @[DCache.scala 49:26]
    end else if (5'h1e == index_addr) begin // @[DCache.scala 120:26]
      v1_30 <= _d1_T | _GEN_67; // @[DCache.scala 120:26]
    end
    if (reset) begin // @[DCache.scala 49:26]
      v1_31 <= 1'h0; // @[DCache.scala 49:26]
    end else if (5'h1f == index_addr) begin // @[DCache.scala 120:26]
      v1_31 <= _d1_T | _GEN_67; // @[DCache.scala 120:26]
    end
    if (reset) begin // @[DCache.scala 50:26]
      d1_0 <= 1'h0; // @[DCache.scala 50:26]
    end else if (5'h0 == index_addr) begin // @[DCache.scala 106:20]
      if (update & updateway1) begin // @[DCache.scala 106:26]
        d1_0 <= 1'h0;
      end else begin
        d1_0 <= way1write | _GEN_355;
      end
    end
    if (reset) begin // @[DCache.scala 50:26]
      d1_1 <= 1'h0; // @[DCache.scala 50:26]
    end else if (5'h1 == index_addr) begin // @[DCache.scala 106:20]
      if (update & updateway1) begin // @[DCache.scala 106:26]
        d1_1 <= 1'h0;
      end else begin
        d1_1 <= way1write | _GEN_355;
      end
    end
    if (reset) begin // @[DCache.scala 50:26]
      d1_2 <= 1'h0; // @[DCache.scala 50:26]
    end else if (5'h2 == index_addr) begin // @[DCache.scala 106:20]
      if (update & updateway1) begin // @[DCache.scala 106:26]
        d1_2 <= 1'h0;
      end else begin
        d1_2 <= way1write | _GEN_355;
      end
    end
    if (reset) begin // @[DCache.scala 50:26]
      d1_3 <= 1'h0; // @[DCache.scala 50:26]
    end else if (5'h3 == index_addr) begin // @[DCache.scala 106:20]
      if (update & updateway1) begin // @[DCache.scala 106:26]
        d1_3 <= 1'h0;
      end else begin
        d1_3 <= way1write | _GEN_355;
      end
    end
    if (reset) begin // @[DCache.scala 50:26]
      d1_4 <= 1'h0; // @[DCache.scala 50:26]
    end else if (5'h4 == index_addr) begin // @[DCache.scala 106:20]
      if (update & updateway1) begin // @[DCache.scala 106:26]
        d1_4 <= 1'h0;
      end else begin
        d1_4 <= way1write | _GEN_355;
      end
    end
    if (reset) begin // @[DCache.scala 50:26]
      d1_5 <= 1'h0; // @[DCache.scala 50:26]
    end else if (5'h5 == index_addr) begin // @[DCache.scala 106:20]
      if (update & updateway1) begin // @[DCache.scala 106:26]
        d1_5 <= 1'h0;
      end else begin
        d1_5 <= way1write | _GEN_355;
      end
    end
    if (reset) begin // @[DCache.scala 50:26]
      d1_6 <= 1'h0; // @[DCache.scala 50:26]
    end else if (5'h6 == index_addr) begin // @[DCache.scala 106:20]
      if (update & updateway1) begin // @[DCache.scala 106:26]
        d1_6 <= 1'h0;
      end else begin
        d1_6 <= way1write | _GEN_355;
      end
    end
    if (reset) begin // @[DCache.scala 50:26]
      d1_7 <= 1'h0; // @[DCache.scala 50:26]
    end else if (5'h7 == index_addr) begin // @[DCache.scala 106:20]
      if (update & updateway1) begin // @[DCache.scala 106:26]
        d1_7 <= 1'h0;
      end else begin
        d1_7 <= way1write | _GEN_355;
      end
    end
    if (reset) begin // @[DCache.scala 50:26]
      d1_8 <= 1'h0; // @[DCache.scala 50:26]
    end else if (5'h8 == index_addr) begin // @[DCache.scala 106:20]
      if (update & updateway1) begin // @[DCache.scala 106:26]
        d1_8 <= 1'h0;
      end else begin
        d1_8 <= way1write | _GEN_355;
      end
    end
    if (reset) begin // @[DCache.scala 50:26]
      d1_9 <= 1'h0; // @[DCache.scala 50:26]
    end else if (5'h9 == index_addr) begin // @[DCache.scala 106:20]
      if (update & updateway1) begin // @[DCache.scala 106:26]
        d1_9 <= 1'h0;
      end else begin
        d1_9 <= way1write | _GEN_355;
      end
    end
    if (reset) begin // @[DCache.scala 50:26]
      d1_10 <= 1'h0; // @[DCache.scala 50:26]
    end else if (5'ha == index_addr) begin // @[DCache.scala 106:20]
      if (update & updateway1) begin // @[DCache.scala 106:26]
        d1_10 <= 1'h0;
      end else begin
        d1_10 <= way1write | _GEN_355;
      end
    end
    if (reset) begin // @[DCache.scala 50:26]
      d1_11 <= 1'h0; // @[DCache.scala 50:26]
    end else if (5'hb == index_addr) begin // @[DCache.scala 106:20]
      if (update & updateway1) begin // @[DCache.scala 106:26]
        d1_11 <= 1'h0;
      end else begin
        d1_11 <= way1write | _GEN_355;
      end
    end
    if (reset) begin // @[DCache.scala 50:26]
      d1_12 <= 1'h0; // @[DCache.scala 50:26]
    end else if (5'hc == index_addr) begin // @[DCache.scala 106:20]
      if (update & updateway1) begin // @[DCache.scala 106:26]
        d1_12 <= 1'h0;
      end else begin
        d1_12 <= way1write | _GEN_355;
      end
    end
    if (reset) begin // @[DCache.scala 50:26]
      d1_13 <= 1'h0; // @[DCache.scala 50:26]
    end else if (5'hd == index_addr) begin // @[DCache.scala 106:20]
      if (update & updateway1) begin // @[DCache.scala 106:26]
        d1_13 <= 1'h0;
      end else begin
        d1_13 <= way1write | _GEN_355;
      end
    end
    if (reset) begin // @[DCache.scala 50:26]
      d1_14 <= 1'h0; // @[DCache.scala 50:26]
    end else if (5'he == index_addr) begin // @[DCache.scala 106:20]
      if (update & updateway1) begin // @[DCache.scala 106:26]
        d1_14 <= 1'h0;
      end else begin
        d1_14 <= way1write | _GEN_355;
      end
    end
    if (reset) begin // @[DCache.scala 50:26]
      d1_15 <= 1'h0; // @[DCache.scala 50:26]
    end else if (5'hf == index_addr) begin // @[DCache.scala 106:20]
      if (update & updateway1) begin // @[DCache.scala 106:26]
        d1_15 <= 1'h0;
      end else begin
        d1_15 <= way1write | _GEN_355;
      end
    end
    if (reset) begin // @[DCache.scala 50:26]
      d1_16 <= 1'h0; // @[DCache.scala 50:26]
    end else if (5'h10 == index_addr) begin // @[DCache.scala 106:20]
      if (update & updateway1) begin // @[DCache.scala 106:26]
        d1_16 <= 1'h0;
      end else begin
        d1_16 <= way1write | _GEN_355;
      end
    end
    if (reset) begin // @[DCache.scala 50:26]
      d1_17 <= 1'h0; // @[DCache.scala 50:26]
    end else if (5'h11 == index_addr) begin // @[DCache.scala 106:20]
      if (update & updateway1) begin // @[DCache.scala 106:26]
        d1_17 <= 1'h0;
      end else begin
        d1_17 <= way1write | _GEN_355;
      end
    end
    if (reset) begin // @[DCache.scala 50:26]
      d1_18 <= 1'h0; // @[DCache.scala 50:26]
    end else if (5'h12 == index_addr) begin // @[DCache.scala 106:20]
      if (update & updateway1) begin // @[DCache.scala 106:26]
        d1_18 <= 1'h0;
      end else begin
        d1_18 <= way1write | _GEN_355;
      end
    end
    if (reset) begin // @[DCache.scala 50:26]
      d1_19 <= 1'h0; // @[DCache.scala 50:26]
    end else if (5'h13 == index_addr) begin // @[DCache.scala 106:20]
      if (update & updateway1) begin // @[DCache.scala 106:26]
        d1_19 <= 1'h0;
      end else begin
        d1_19 <= way1write | _GEN_355;
      end
    end
    if (reset) begin // @[DCache.scala 50:26]
      d1_20 <= 1'h0; // @[DCache.scala 50:26]
    end else if (5'h14 == index_addr) begin // @[DCache.scala 106:20]
      if (update & updateway1) begin // @[DCache.scala 106:26]
        d1_20 <= 1'h0;
      end else begin
        d1_20 <= way1write | _GEN_355;
      end
    end
    if (reset) begin // @[DCache.scala 50:26]
      d1_21 <= 1'h0; // @[DCache.scala 50:26]
    end else if (5'h15 == index_addr) begin // @[DCache.scala 106:20]
      if (update & updateway1) begin // @[DCache.scala 106:26]
        d1_21 <= 1'h0;
      end else begin
        d1_21 <= way1write | _GEN_355;
      end
    end
    if (reset) begin // @[DCache.scala 50:26]
      d1_22 <= 1'h0; // @[DCache.scala 50:26]
    end else if (5'h16 == index_addr) begin // @[DCache.scala 106:20]
      if (update & updateway1) begin // @[DCache.scala 106:26]
        d1_22 <= 1'h0;
      end else begin
        d1_22 <= way1write | _GEN_355;
      end
    end
    if (reset) begin // @[DCache.scala 50:26]
      d1_23 <= 1'h0; // @[DCache.scala 50:26]
    end else if (5'h17 == index_addr) begin // @[DCache.scala 106:20]
      if (update & updateway1) begin // @[DCache.scala 106:26]
        d1_23 <= 1'h0;
      end else begin
        d1_23 <= way1write | _GEN_355;
      end
    end
    if (reset) begin // @[DCache.scala 50:26]
      d1_24 <= 1'h0; // @[DCache.scala 50:26]
    end else if (5'h18 == index_addr) begin // @[DCache.scala 106:20]
      if (update & updateway1) begin // @[DCache.scala 106:26]
        d1_24 <= 1'h0;
      end else begin
        d1_24 <= way1write | _GEN_355;
      end
    end
    if (reset) begin // @[DCache.scala 50:26]
      d1_25 <= 1'h0; // @[DCache.scala 50:26]
    end else if (5'h19 == index_addr) begin // @[DCache.scala 106:20]
      if (update & updateway1) begin // @[DCache.scala 106:26]
        d1_25 <= 1'h0;
      end else begin
        d1_25 <= way1write | _GEN_355;
      end
    end
    if (reset) begin // @[DCache.scala 50:26]
      d1_26 <= 1'h0; // @[DCache.scala 50:26]
    end else if (5'h1a == index_addr) begin // @[DCache.scala 106:20]
      if (update & updateway1) begin // @[DCache.scala 106:26]
        d1_26 <= 1'h0;
      end else begin
        d1_26 <= way1write | _GEN_355;
      end
    end
    if (reset) begin // @[DCache.scala 50:26]
      d1_27 <= 1'h0; // @[DCache.scala 50:26]
    end else if (5'h1b == index_addr) begin // @[DCache.scala 106:20]
      if (update & updateway1) begin // @[DCache.scala 106:26]
        d1_27 <= 1'h0;
      end else begin
        d1_27 <= way1write | _GEN_355;
      end
    end
    if (reset) begin // @[DCache.scala 50:26]
      d1_28 <= 1'h0; // @[DCache.scala 50:26]
    end else if (5'h1c == index_addr) begin // @[DCache.scala 106:20]
      if (update & updateway1) begin // @[DCache.scala 106:26]
        d1_28 <= 1'h0;
      end else begin
        d1_28 <= way1write | _GEN_355;
      end
    end
    if (reset) begin // @[DCache.scala 50:26]
      d1_29 <= 1'h0; // @[DCache.scala 50:26]
    end else if (5'h1d == index_addr) begin // @[DCache.scala 106:20]
      if (update & updateway1) begin // @[DCache.scala 106:26]
        d1_29 <= 1'h0;
      end else begin
        d1_29 <= way1write | _GEN_355;
      end
    end
    if (reset) begin // @[DCache.scala 50:26]
      d1_30 <= 1'h0; // @[DCache.scala 50:26]
    end else if (5'h1e == index_addr) begin // @[DCache.scala 106:20]
      if (update & updateway1) begin // @[DCache.scala 106:26]
        d1_30 <= 1'h0;
      end else begin
        d1_30 <= way1write | _GEN_355;
      end
    end
    if (reset) begin // @[DCache.scala 50:26]
      d1_31 <= 1'h0; // @[DCache.scala 50:26]
    end else if (5'h1f == index_addr) begin // @[DCache.scala 106:20]
      if (update & updateway1) begin // @[DCache.scala 106:26]
        d1_31 <= 1'h0;
      end else begin
        d1_31 <= way1write | _GEN_355;
      end
    end
    if (reset) begin // @[DCache.scala 51:26]
      age1_0 <= 1'h0; // @[DCache.scala 51:26]
    end else if (5'h0 == index_addr) begin // @[DCache.scala 78:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 78:28]
        age1_0 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 78:28]
        age1_0 <= age1_31; // @[DCache.scala 78:28]
      end else begin
        age1_0 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 51:26]
      age1_1 <= 1'h0; // @[DCache.scala 51:26]
    end else if (5'h1 == index_addr) begin // @[DCache.scala 78:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 78:28]
        age1_1 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 78:28]
        age1_1 <= age1_31; // @[DCache.scala 78:28]
      end else begin
        age1_1 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 51:26]
      age1_2 <= 1'h0; // @[DCache.scala 51:26]
    end else if (5'h2 == index_addr) begin // @[DCache.scala 78:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 78:28]
        age1_2 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 78:28]
        age1_2 <= age1_31; // @[DCache.scala 78:28]
      end else begin
        age1_2 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 51:26]
      age1_3 <= 1'h0; // @[DCache.scala 51:26]
    end else if (5'h3 == index_addr) begin // @[DCache.scala 78:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 78:28]
        age1_3 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 78:28]
        age1_3 <= age1_31; // @[DCache.scala 78:28]
      end else begin
        age1_3 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 51:26]
      age1_4 <= 1'h0; // @[DCache.scala 51:26]
    end else if (5'h4 == index_addr) begin // @[DCache.scala 78:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 78:28]
        age1_4 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 78:28]
        age1_4 <= age1_31; // @[DCache.scala 78:28]
      end else begin
        age1_4 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 51:26]
      age1_5 <= 1'h0; // @[DCache.scala 51:26]
    end else if (5'h5 == index_addr) begin // @[DCache.scala 78:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 78:28]
        age1_5 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 78:28]
        age1_5 <= age1_31; // @[DCache.scala 78:28]
      end else begin
        age1_5 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 51:26]
      age1_6 <= 1'h0; // @[DCache.scala 51:26]
    end else if (5'h6 == index_addr) begin // @[DCache.scala 78:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 78:28]
        age1_6 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 78:28]
        age1_6 <= age1_31; // @[DCache.scala 78:28]
      end else begin
        age1_6 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 51:26]
      age1_7 <= 1'h0; // @[DCache.scala 51:26]
    end else if (5'h7 == index_addr) begin // @[DCache.scala 78:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 78:28]
        age1_7 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 78:28]
        age1_7 <= age1_31; // @[DCache.scala 78:28]
      end else begin
        age1_7 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 51:26]
      age1_8 <= 1'h0; // @[DCache.scala 51:26]
    end else if (5'h8 == index_addr) begin // @[DCache.scala 78:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 78:28]
        age1_8 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 78:28]
        age1_8 <= age1_31; // @[DCache.scala 78:28]
      end else begin
        age1_8 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 51:26]
      age1_9 <= 1'h0; // @[DCache.scala 51:26]
    end else if (5'h9 == index_addr) begin // @[DCache.scala 78:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 78:28]
        age1_9 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 78:28]
        age1_9 <= age1_31; // @[DCache.scala 78:28]
      end else begin
        age1_9 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 51:26]
      age1_10 <= 1'h0; // @[DCache.scala 51:26]
    end else if (5'ha == index_addr) begin // @[DCache.scala 78:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 78:28]
        age1_10 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 78:28]
        age1_10 <= age1_31; // @[DCache.scala 78:28]
      end else begin
        age1_10 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 51:26]
      age1_11 <= 1'h0; // @[DCache.scala 51:26]
    end else if (5'hb == index_addr) begin // @[DCache.scala 78:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 78:28]
        age1_11 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 78:28]
        age1_11 <= age1_31; // @[DCache.scala 78:28]
      end else begin
        age1_11 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 51:26]
      age1_12 <= 1'h0; // @[DCache.scala 51:26]
    end else if (5'hc == index_addr) begin // @[DCache.scala 78:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 78:28]
        age1_12 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 78:28]
        age1_12 <= age1_31; // @[DCache.scala 78:28]
      end else begin
        age1_12 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 51:26]
      age1_13 <= 1'h0; // @[DCache.scala 51:26]
    end else if (5'hd == index_addr) begin // @[DCache.scala 78:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 78:28]
        age1_13 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 78:28]
        age1_13 <= age1_31; // @[DCache.scala 78:28]
      end else begin
        age1_13 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 51:26]
      age1_14 <= 1'h0; // @[DCache.scala 51:26]
    end else if (5'he == index_addr) begin // @[DCache.scala 78:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 78:28]
        age1_14 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 78:28]
        age1_14 <= age1_31; // @[DCache.scala 78:28]
      end else begin
        age1_14 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 51:26]
      age1_15 <= 1'h0; // @[DCache.scala 51:26]
    end else if (5'hf == index_addr) begin // @[DCache.scala 78:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 78:28]
        age1_15 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 78:28]
        age1_15 <= age1_31; // @[DCache.scala 78:28]
      end else begin
        age1_15 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 51:26]
      age1_16 <= 1'h0; // @[DCache.scala 51:26]
    end else if (5'h10 == index_addr) begin // @[DCache.scala 78:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 78:28]
        age1_16 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 78:28]
        age1_16 <= age1_31; // @[DCache.scala 78:28]
      end else begin
        age1_16 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 51:26]
      age1_17 <= 1'h0; // @[DCache.scala 51:26]
    end else if (5'h11 == index_addr) begin // @[DCache.scala 78:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 78:28]
        age1_17 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 78:28]
        age1_17 <= age1_31; // @[DCache.scala 78:28]
      end else begin
        age1_17 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 51:26]
      age1_18 <= 1'h0; // @[DCache.scala 51:26]
    end else if (5'h12 == index_addr) begin // @[DCache.scala 78:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 78:28]
        age1_18 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 78:28]
        age1_18 <= age1_31; // @[DCache.scala 78:28]
      end else begin
        age1_18 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 51:26]
      age1_19 <= 1'h0; // @[DCache.scala 51:26]
    end else if (5'h13 == index_addr) begin // @[DCache.scala 78:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 78:28]
        age1_19 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 78:28]
        age1_19 <= age1_31; // @[DCache.scala 78:28]
      end else begin
        age1_19 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 51:26]
      age1_20 <= 1'h0; // @[DCache.scala 51:26]
    end else if (5'h14 == index_addr) begin // @[DCache.scala 78:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 78:28]
        age1_20 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 78:28]
        age1_20 <= age1_31; // @[DCache.scala 78:28]
      end else begin
        age1_20 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 51:26]
      age1_21 <= 1'h0; // @[DCache.scala 51:26]
    end else if (5'h15 == index_addr) begin // @[DCache.scala 78:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 78:28]
        age1_21 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 78:28]
        age1_21 <= age1_31; // @[DCache.scala 78:28]
      end else begin
        age1_21 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 51:26]
      age1_22 <= 1'h0; // @[DCache.scala 51:26]
    end else if (5'h16 == index_addr) begin // @[DCache.scala 78:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 78:28]
        age1_22 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 78:28]
        age1_22 <= age1_31; // @[DCache.scala 78:28]
      end else begin
        age1_22 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 51:26]
      age1_23 <= 1'h0; // @[DCache.scala 51:26]
    end else if (5'h17 == index_addr) begin // @[DCache.scala 78:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 78:28]
        age1_23 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 78:28]
        age1_23 <= age1_31; // @[DCache.scala 78:28]
      end else begin
        age1_23 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 51:26]
      age1_24 <= 1'h0; // @[DCache.scala 51:26]
    end else if (5'h18 == index_addr) begin // @[DCache.scala 78:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 78:28]
        age1_24 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 78:28]
        age1_24 <= age1_31; // @[DCache.scala 78:28]
      end else begin
        age1_24 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 51:26]
      age1_25 <= 1'h0; // @[DCache.scala 51:26]
    end else if (5'h19 == index_addr) begin // @[DCache.scala 78:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 78:28]
        age1_25 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 78:28]
        age1_25 <= age1_31; // @[DCache.scala 78:28]
      end else begin
        age1_25 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 51:26]
      age1_26 <= 1'h0; // @[DCache.scala 51:26]
    end else if (5'h1a == index_addr) begin // @[DCache.scala 78:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 78:28]
        age1_26 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 78:28]
        age1_26 <= age1_31; // @[DCache.scala 78:28]
      end else begin
        age1_26 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 51:26]
      age1_27 <= 1'h0; // @[DCache.scala 51:26]
    end else if (5'h1b == index_addr) begin // @[DCache.scala 78:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 78:28]
        age1_27 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 78:28]
        age1_27 <= age1_31; // @[DCache.scala 78:28]
      end else begin
        age1_27 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 51:26]
      age1_28 <= 1'h0; // @[DCache.scala 51:26]
    end else if (5'h1c == index_addr) begin // @[DCache.scala 78:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 78:28]
        age1_28 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 78:28]
        age1_28 <= age1_31; // @[DCache.scala 78:28]
      end else begin
        age1_28 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 51:26]
      age1_29 <= 1'h0; // @[DCache.scala 51:26]
    end else if (5'h1d == index_addr) begin // @[DCache.scala 78:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 78:28]
        age1_29 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 78:28]
        age1_29 <= age1_31; // @[DCache.scala 78:28]
      end else begin
        age1_29 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 51:26]
      age1_30 <= 1'h0; // @[DCache.scala 51:26]
    end else if (5'h1e == index_addr) begin // @[DCache.scala 78:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 78:28]
        age1_30 <= hit1;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 78:28]
        age1_30 <= age1_31; // @[DCache.scala 78:28]
      end else begin
        age1_30 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 51:26]
      age1_31 <= 1'h0; // @[DCache.scala 51:26]
    end else if (5'h1f == index_addr) begin // @[DCache.scala 78:22]
      if (hit1 ^ hit2) begin // @[DCache.scala 78:28]
        age1_31 <= hit1;
      end else if (!(5'h1f == index_addr)) begin // @[DCache.scala 78:28]
        age1_31 <= _GEN_226;
      end
    end
    if (reset) begin // @[DCache.scala 52:26]
      tag1_0 <= 53'h0; // @[DCache.scala 52:26]
    end else if (5'h0 == index_addr) begin // @[DCache.scala 119:26]
      if (_d1_T) begin // @[DCache.scala 119:32]
        tag1_0 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 60:28]
        tag1_0 <= tag1_31; // @[DCache.scala 60:28]
      end else begin
        tag1_0 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 52:26]
      tag1_1 <= 53'h0; // @[DCache.scala 52:26]
    end else if (5'h1 == index_addr) begin // @[DCache.scala 119:26]
      if (_d1_T) begin // @[DCache.scala 119:32]
        tag1_1 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 60:28]
        tag1_1 <= tag1_31; // @[DCache.scala 60:28]
      end else begin
        tag1_1 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 52:26]
      tag1_2 <= 53'h0; // @[DCache.scala 52:26]
    end else if (5'h2 == index_addr) begin // @[DCache.scala 119:26]
      if (_d1_T) begin // @[DCache.scala 119:32]
        tag1_2 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 60:28]
        tag1_2 <= tag1_31; // @[DCache.scala 60:28]
      end else begin
        tag1_2 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 52:26]
      tag1_3 <= 53'h0; // @[DCache.scala 52:26]
    end else if (5'h3 == index_addr) begin // @[DCache.scala 119:26]
      if (_d1_T) begin // @[DCache.scala 119:32]
        tag1_3 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 60:28]
        tag1_3 <= tag1_31; // @[DCache.scala 60:28]
      end else begin
        tag1_3 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 52:26]
      tag1_4 <= 53'h0; // @[DCache.scala 52:26]
    end else if (5'h4 == index_addr) begin // @[DCache.scala 119:26]
      if (_d1_T) begin // @[DCache.scala 119:32]
        tag1_4 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 60:28]
        tag1_4 <= tag1_31; // @[DCache.scala 60:28]
      end else begin
        tag1_4 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 52:26]
      tag1_5 <= 53'h0; // @[DCache.scala 52:26]
    end else if (5'h5 == index_addr) begin // @[DCache.scala 119:26]
      if (_d1_T) begin // @[DCache.scala 119:32]
        tag1_5 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 60:28]
        tag1_5 <= tag1_31; // @[DCache.scala 60:28]
      end else begin
        tag1_5 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 52:26]
      tag1_6 <= 53'h0; // @[DCache.scala 52:26]
    end else if (5'h6 == index_addr) begin // @[DCache.scala 119:26]
      if (_d1_T) begin // @[DCache.scala 119:32]
        tag1_6 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 60:28]
        tag1_6 <= tag1_31; // @[DCache.scala 60:28]
      end else begin
        tag1_6 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 52:26]
      tag1_7 <= 53'h0; // @[DCache.scala 52:26]
    end else if (5'h7 == index_addr) begin // @[DCache.scala 119:26]
      if (_d1_T) begin // @[DCache.scala 119:32]
        tag1_7 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 60:28]
        tag1_7 <= tag1_31; // @[DCache.scala 60:28]
      end else begin
        tag1_7 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 52:26]
      tag1_8 <= 53'h0; // @[DCache.scala 52:26]
    end else if (5'h8 == index_addr) begin // @[DCache.scala 119:26]
      if (_d1_T) begin // @[DCache.scala 119:32]
        tag1_8 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 60:28]
        tag1_8 <= tag1_31; // @[DCache.scala 60:28]
      end else begin
        tag1_8 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 52:26]
      tag1_9 <= 53'h0; // @[DCache.scala 52:26]
    end else if (5'h9 == index_addr) begin // @[DCache.scala 119:26]
      if (_d1_T) begin // @[DCache.scala 119:32]
        tag1_9 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 60:28]
        tag1_9 <= tag1_31; // @[DCache.scala 60:28]
      end else begin
        tag1_9 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 52:26]
      tag1_10 <= 53'h0; // @[DCache.scala 52:26]
    end else if (5'ha == index_addr) begin // @[DCache.scala 119:26]
      if (_d1_T) begin // @[DCache.scala 119:32]
        tag1_10 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 60:28]
        tag1_10 <= tag1_31; // @[DCache.scala 60:28]
      end else begin
        tag1_10 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 52:26]
      tag1_11 <= 53'h0; // @[DCache.scala 52:26]
    end else if (5'hb == index_addr) begin // @[DCache.scala 119:26]
      if (_d1_T) begin // @[DCache.scala 119:32]
        tag1_11 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 60:28]
        tag1_11 <= tag1_31; // @[DCache.scala 60:28]
      end else begin
        tag1_11 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 52:26]
      tag1_12 <= 53'h0; // @[DCache.scala 52:26]
    end else if (5'hc == index_addr) begin // @[DCache.scala 119:26]
      if (_d1_T) begin // @[DCache.scala 119:32]
        tag1_12 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 60:28]
        tag1_12 <= tag1_31; // @[DCache.scala 60:28]
      end else begin
        tag1_12 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 52:26]
      tag1_13 <= 53'h0; // @[DCache.scala 52:26]
    end else if (5'hd == index_addr) begin // @[DCache.scala 119:26]
      if (_d1_T) begin // @[DCache.scala 119:32]
        tag1_13 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 60:28]
        tag1_13 <= tag1_31; // @[DCache.scala 60:28]
      end else begin
        tag1_13 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 52:26]
      tag1_14 <= 53'h0; // @[DCache.scala 52:26]
    end else if (5'he == index_addr) begin // @[DCache.scala 119:26]
      if (_d1_T) begin // @[DCache.scala 119:32]
        tag1_14 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 60:28]
        tag1_14 <= tag1_31; // @[DCache.scala 60:28]
      end else begin
        tag1_14 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 52:26]
      tag1_15 <= 53'h0; // @[DCache.scala 52:26]
    end else if (5'hf == index_addr) begin // @[DCache.scala 119:26]
      if (_d1_T) begin // @[DCache.scala 119:32]
        tag1_15 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 60:28]
        tag1_15 <= tag1_31; // @[DCache.scala 60:28]
      end else begin
        tag1_15 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 52:26]
      tag1_16 <= 53'h0; // @[DCache.scala 52:26]
    end else if (5'h10 == index_addr) begin // @[DCache.scala 119:26]
      if (_d1_T) begin // @[DCache.scala 119:32]
        tag1_16 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 60:28]
        tag1_16 <= tag1_31; // @[DCache.scala 60:28]
      end else begin
        tag1_16 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 52:26]
      tag1_17 <= 53'h0; // @[DCache.scala 52:26]
    end else if (5'h11 == index_addr) begin // @[DCache.scala 119:26]
      if (_d1_T) begin // @[DCache.scala 119:32]
        tag1_17 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 60:28]
        tag1_17 <= tag1_31; // @[DCache.scala 60:28]
      end else begin
        tag1_17 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 52:26]
      tag1_18 <= 53'h0; // @[DCache.scala 52:26]
    end else if (5'h12 == index_addr) begin // @[DCache.scala 119:26]
      if (_d1_T) begin // @[DCache.scala 119:32]
        tag1_18 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 60:28]
        tag1_18 <= tag1_31; // @[DCache.scala 60:28]
      end else begin
        tag1_18 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 52:26]
      tag1_19 <= 53'h0; // @[DCache.scala 52:26]
    end else if (5'h13 == index_addr) begin // @[DCache.scala 119:26]
      if (_d1_T) begin // @[DCache.scala 119:32]
        tag1_19 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 60:28]
        tag1_19 <= tag1_31; // @[DCache.scala 60:28]
      end else begin
        tag1_19 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 52:26]
      tag1_20 <= 53'h0; // @[DCache.scala 52:26]
    end else if (5'h14 == index_addr) begin // @[DCache.scala 119:26]
      if (_d1_T) begin // @[DCache.scala 119:32]
        tag1_20 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 60:28]
        tag1_20 <= tag1_31; // @[DCache.scala 60:28]
      end else begin
        tag1_20 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 52:26]
      tag1_21 <= 53'h0; // @[DCache.scala 52:26]
    end else if (5'h15 == index_addr) begin // @[DCache.scala 119:26]
      if (_d1_T) begin // @[DCache.scala 119:32]
        tag1_21 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 60:28]
        tag1_21 <= tag1_31; // @[DCache.scala 60:28]
      end else begin
        tag1_21 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 52:26]
      tag1_22 <= 53'h0; // @[DCache.scala 52:26]
    end else if (5'h16 == index_addr) begin // @[DCache.scala 119:26]
      if (_d1_T) begin // @[DCache.scala 119:32]
        tag1_22 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 60:28]
        tag1_22 <= tag1_31; // @[DCache.scala 60:28]
      end else begin
        tag1_22 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 52:26]
      tag1_23 <= 53'h0; // @[DCache.scala 52:26]
    end else if (5'h17 == index_addr) begin // @[DCache.scala 119:26]
      if (_d1_T) begin // @[DCache.scala 119:32]
        tag1_23 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 60:28]
        tag1_23 <= tag1_31; // @[DCache.scala 60:28]
      end else begin
        tag1_23 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 52:26]
      tag1_24 <= 53'h0; // @[DCache.scala 52:26]
    end else if (5'h18 == index_addr) begin // @[DCache.scala 119:26]
      if (_d1_T) begin // @[DCache.scala 119:32]
        tag1_24 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 60:28]
        tag1_24 <= tag1_31; // @[DCache.scala 60:28]
      end else begin
        tag1_24 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 52:26]
      tag1_25 <= 53'h0; // @[DCache.scala 52:26]
    end else if (5'h19 == index_addr) begin // @[DCache.scala 119:26]
      if (_d1_T) begin // @[DCache.scala 119:32]
        tag1_25 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 60:28]
        tag1_25 <= tag1_31; // @[DCache.scala 60:28]
      end else begin
        tag1_25 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 52:26]
      tag1_26 <= 53'h0; // @[DCache.scala 52:26]
    end else if (5'h1a == index_addr) begin // @[DCache.scala 119:26]
      if (_d1_T) begin // @[DCache.scala 119:32]
        tag1_26 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 60:28]
        tag1_26 <= tag1_31; // @[DCache.scala 60:28]
      end else begin
        tag1_26 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 52:26]
      tag1_27 <= 53'h0; // @[DCache.scala 52:26]
    end else if (5'h1b == index_addr) begin // @[DCache.scala 119:26]
      if (_d1_T) begin // @[DCache.scala 119:32]
        tag1_27 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 60:28]
        tag1_27 <= tag1_31; // @[DCache.scala 60:28]
      end else begin
        tag1_27 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 52:26]
      tag1_28 <= 53'h0; // @[DCache.scala 52:26]
    end else if (5'h1c == index_addr) begin // @[DCache.scala 119:26]
      if (_d1_T) begin // @[DCache.scala 119:32]
        tag1_28 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 60:28]
        tag1_28 <= tag1_31; // @[DCache.scala 60:28]
      end else begin
        tag1_28 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 52:26]
      tag1_29 <= 53'h0; // @[DCache.scala 52:26]
    end else if (5'h1d == index_addr) begin // @[DCache.scala 119:26]
      if (_d1_T) begin // @[DCache.scala 119:32]
        tag1_29 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 60:28]
        tag1_29 <= tag1_31; // @[DCache.scala 60:28]
      end else begin
        tag1_29 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 52:26]
      tag1_30 <= 53'h0; // @[DCache.scala 52:26]
    end else if (5'h1e == index_addr) begin // @[DCache.scala 119:26]
      if (_d1_T) begin // @[DCache.scala 119:32]
        tag1_30 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 60:28]
        tag1_30 <= tag1_31; // @[DCache.scala 60:28]
      end else begin
        tag1_30 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 52:26]
      tag1_31 <= 53'h0; // @[DCache.scala 52:26]
    end else if (5'h1f == index_addr) begin // @[DCache.scala 119:26]
      if (_d1_T) begin // @[DCache.scala 119:32]
        tag1_31 <= tag_addr;
      end else if (!(5'h1f == index_addr)) begin // @[DCache.scala 60:28]
        tag1_31 <= _GEN_34;
      end
    end
    if (reset) begin // @[DCache.scala 53:26]
      block1_0 <= 512'h0; // @[DCache.scala 53:26]
    end else if (5'h0 == index_addr) begin // @[DCache.scala 118:26]
      if (_d1_T) begin // @[DCache.scala 118:32]
        block1_0 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 118:72]
        block1_0 <= block1_after_write;
      end else begin
        block1_0 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 53:26]
      block1_1 <= 512'h0; // @[DCache.scala 53:26]
    end else if (5'h1 == index_addr) begin // @[DCache.scala 118:26]
      if (_d1_T) begin // @[DCache.scala 118:32]
        block1_1 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 118:72]
        block1_1 <= block1_after_write;
      end else begin
        block1_1 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 53:26]
      block1_2 <= 512'h0; // @[DCache.scala 53:26]
    end else if (5'h2 == index_addr) begin // @[DCache.scala 118:26]
      if (_d1_T) begin // @[DCache.scala 118:32]
        block1_2 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 118:72]
        block1_2 <= block1_after_write;
      end else begin
        block1_2 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 53:26]
      block1_3 <= 512'h0; // @[DCache.scala 53:26]
    end else if (5'h3 == index_addr) begin // @[DCache.scala 118:26]
      if (_d1_T) begin // @[DCache.scala 118:32]
        block1_3 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 118:72]
        block1_3 <= block1_after_write;
      end else begin
        block1_3 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 53:26]
      block1_4 <= 512'h0; // @[DCache.scala 53:26]
    end else if (5'h4 == index_addr) begin // @[DCache.scala 118:26]
      if (_d1_T) begin // @[DCache.scala 118:32]
        block1_4 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 118:72]
        block1_4 <= block1_after_write;
      end else begin
        block1_4 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 53:26]
      block1_5 <= 512'h0; // @[DCache.scala 53:26]
    end else if (5'h5 == index_addr) begin // @[DCache.scala 118:26]
      if (_d1_T) begin // @[DCache.scala 118:32]
        block1_5 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 118:72]
        block1_5 <= block1_after_write;
      end else begin
        block1_5 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 53:26]
      block1_6 <= 512'h0; // @[DCache.scala 53:26]
    end else if (5'h6 == index_addr) begin // @[DCache.scala 118:26]
      if (_d1_T) begin // @[DCache.scala 118:32]
        block1_6 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 118:72]
        block1_6 <= block1_after_write;
      end else begin
        block1_6 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 53:26]
      block1_7 <= 512'h0; // @[DCache.scala 53:26]
    end else if (5'h7 == index_addr) begin // @[DCache.scala 118:26]
      if (_d1_T) begin // @[DCache.scala 118:32]
        block1_7 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 118:72]
        block1_7 <= block1_after_write;
      end else begin
        block1_7 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 53:26]
      block1_8 <= 512'h0; // @[DCache.scala 53:26]
    end else if (5'h8 == index_addr) begin // @[DCache.scala 118:26]
      if (_d1_T) begin // @[DCache.scala 118:32]
        block1_8 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 118:72]
        block1_8 <= block1_after_write;
      end else begin
        block1_8 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 53:26]
      block1_9 <= 512'h0; // @[DCache.scala 53:26]
    end else if (5'h9 == index_addr) begin // @[DCache.scala 118:26]
      if (_d1_T) begin // @[DCache.scala 118:32]
        block1_9 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 118:72]
        block1_9 <= block1_after_write;
      end else begin
        block1_9 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 53:26]
      block1_10 <= 512'h0; // @[DCache.scala 53:26]
    end else if (5'ha == index_addr) begin // @[DCache.scala 118:26]
      if (_d1_T) begin // @[DCache.scala 118:32]
        block1_10 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 118:72]
        block1_10 <= block1_after_write;
      end else begin
        block1_10 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 53:26]
      block1_11 <= 512'h0; // @[DCache.scala 53:26]
    end else if (5'hb == index_addr) begin // @[DCache.scala 118:26]
      if (_d1_T) begin // @[DCache.scala 118:32]
        block1_11 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 118:72]
        block1_11 <= block1_after_write;
      end else begin
        block1_11 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 53:26]
      block1_12 <= 512'h0; // @[DCache.scala 53:26]
    end else if (5'hc == index_addr) begin // @[DCache.scala 118:26]
      if (_d1_T) begin // @[DCache.scala 118:32]
        block1_12 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 118:72]
        block1_12 <= block1_after_write;
      end else begin
        block1_12 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 53:26]
      block1_13 <= 512'h0; // @[DCache.scala 53:26]
    end else if (5'hd == index_addr) begin // @[DCache.scala 118:26]
      if (_d1_T) begin // @[DCache.scala 118:32]
        block1_13 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 118:72]
        block1_13 <= block1_after_write;
      end else begin
        block1_13 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 53:26]
      block1_14 <= 512'h0; // @[DCache.scala 53:26]
    end else if (5'he == index_addr) begin // @[DCache.scala 118:26]
      if (_d1_T) begin // @[DCache.scala 118:32]
        block1_14 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 118:72]
        block1_14 <= block1_after_write;
      end else begin
        block1_14 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 53:26]
      block1_15 <= 512'h0; // @[DCache.scala 53:26]
    end else if (5'hf == index_addr) begin // @[DCache.scala 118:26]
      if (_d1_T) begin // @[DCache.scala 118:32]
        block1_15 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 118:72]
        block1_15 <= block1_after_write;
      end else begin
        block1_15 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 53:26]
      block1_16 <= 512'h0; // @[DCache.scala 53:26]
    end else if (5'h10 == index_addr) begin // @[DCache.scala 118:26]
      if (_d1_T) begin // @[DCache.scala 118:32]
        block1_16 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 118:72]
        block1_16 <= block1_after_write;
      end else begin
        block1_16 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 53:26]
      block1_17 <= 512'h0; // @[DCache.scala 53:26]
    end else if (5'h11 == index_addr) begin // @[DCache.scala 118:26]
      if (_d1_T) begin // @[DCache.scala 118:32]
        block1_17 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 118:72]
        block1_17 <= block1_after_write;
      end else begin
        block1_17 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 53:26]
      block1_18 <= 512'h0; // @[DCache.scala 53:26]
    end else if (5'h12 == index_addr) begin // @[DCache.scala 118:26]
      if (_d1_T) begin // @[DCache.scala 118:32]
        block1_18 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 118:72]
        block1_18 <= block1_after_write;
      end else begin
        block1_18 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 53:26]
      block1_19 <= 512'h0; // @[DCache.scala 53:26]
    end else if (5'h13 == index_addr) begin // @[DCache.scala 118:26]
      if (_d1_T) begin // @[DCache.scala 118:32]
        block1_19 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 118:72]
        block1_19 <= block1_after_write;
      end else begin
        block1_19 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 53:26]
      block1_20 <= 512'h0; // @[DCache.scala 53:26]
    end else if (5'h14 == index_addr) begin // @[DCache.scala 118:26]
      if (_d1_T) begin // @[DCache.scala 118:32]
        block1_20 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 118:72]
        block1_20 <= block1_after_write;
      end else begin
        block1_20 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 53:26]
      block1_21 <= 512'h0; // @[DCache.scala 53:26]
    end else if (5'h15 == index_addr) begin // @[DCache.scala 118:26]
      if (_d1_T) begin // @[DCache.scala 118:32]
        block1_21 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 118:72]
        block1_21 <= block1_after_write;
      end else begin
        block1_21 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 53:26]
      block1_22 <= 512'h0; // @[DCache.scala 53:26]
    end else if (5'h16 == index_addr) begin // @[DCache.scala 118:26]
      if (_d1_T) begin // @[DCache.scala 118:32]
        block1_22 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 118:72]
        block1_22 <= block1_after_write;
      end else begin
        block1_22 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 53:26]
      block1_23 <= 512'h0; // @[DCache.scala 53:26]
    end else if (5'h17 == index_addr) begin // @[DCache.scala 118:26]
      if (_d1_T) begin // @[DCache.scala 118:32]
        block1_23 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 118:72]
        block1_23 <= block1_after_write;
      end else begin
        block1_23 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 53:26]
      block1_24 <= 512'h0; // @[DCache.scala 53:26]
    end else if (5'h18 == index_addr) begin // @[DCache.scala 118:26]
      if (_d1_T) begin // @[DCache.scala 118:32]
        block1_24 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 118:72]
        block1_24 <= block1_after_write;
      end else begin
        block1_24 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 53:26]
      block1_25 <= 512'h0; // @[DCache.scala 53:26]
    end else if (5'h19 == index_addr) begin // @[DCache.scala 118:26]
      if (_d1_T) begin // @[DCache.scala 118:32]
        block1_25 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 118:72]
        block1_25 <= block1_after_write;
      end else begin
        block1_25 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 53:26]
      block1_26 <= 512'h0; // @[DCache.scala 53:26]
    end else if (5'h1a == index_addr) begin // @[DCache.scala 118:26]
      if (_d1_T) begin // @[DCache.scala 118:32]
        block1_26 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 118:72]
        block1_26 <= block1_after_write;
      end else begin
        block1_26 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 53:26]
      block1_27 <= 512'h0; // @[DCache.scala 53:26]
    end else if (5'h1b == index_addr) begin // @[DCache.scala 118:26]
      if (_d1_T) begin // @[DCache.scala 118:32]
        block1_27 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 118:72]
        block1_27 <= block1_after_write;
      end else begin
        block1_27 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 53:26]
      block1_28 <= 512'h0; // @[DCache.scala 53:26]
    end else if (5'h1c == index_addr) begin // @[DCache.scala 118:26]
      if (_d1_T) begin // @[DCache.scala 118:32]
        block1_28 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 118:72]
        block1_28 <= block1_after_write;
      end else begin
        block1_28 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 53:26]
      block1_29 <= 512'h0; // @[DCache.scala 53:26]
    end else if (5'h1d == index_addr) begin // @[DCache.scala 118:26]
      if (_d1_T) begin // @[DCache.scala 118:32]
        block1_29 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 118:72]
        block1_29 <= block1_after_write;
      end else begin
        block1_29 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 53:26]
      block1_30 <= 512'h0; // @[DCache.scala 53:26]
    end else if (5'h1e == index_addr) begin // @[DCache.scala 118:26]
      if (_d1_T) begin // @[DCache.scala 118:32]
        block1_30 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 118:72]
        block1_30 <= block1_after_write;
      end else begin
        block1_30 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 53:26]
      block1_31 <= 512'h0; // @[DCache.scala 53:26]
    end else if (5'h1f == index_addr) begin // @[DCache.scala 118:26]
      if (_d1_T) begin // @[DCache.scala 118:32]
        block1_31 <= io_axi_rdata;
      end else if (way1write) begin // @[DCache.scala 118:72]
        block1_31 <= block1_after_write;
      end else begin
        block1_31 <= _GEN_163;
      end
    end
    if (reset) begin // @[DCache.scala 54:26]
      v2_0 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h0 == index_addr) begin // @[DCache.scala 123:26]
      v2_0 <= _d2_T | _GEN_131; // @[DCache.scala 123:26]
    end
    if (reset) begin // @[DCache.scala 54:26]
      v2_1 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h1 == index_addr) begin // @[DCache.scala 123:26]
      v2_1 <= _d2_T | _GEN_131; // @[DCache.scala 123:26]
    end
    if (reset) begin // @[DCache.scala 54:26]
      v2_2 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h2 == index_addr) begin // @[DCache.scala 123:26]
      v2_2 <= _d2_T | _GEN_131; // @[DCache.scala 123:26]
    end
    if (reset) begin // @[DCache.scala 54:26]
      v2_3 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h3 == index_addr) begin // @[DCache.scala 123:26]
      v2_3 <= _d2_T | _GEN_131; // @[DCache.scala 123:26]
    end
    if (reset) begin // @[DCache.scala 54:26]
      v2_4 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h4 == index_addr) begin // @[DCache.scala 123:26]
      v2_4 <= _d2_T | _GEN_131; // @[DCache.scala 123:26]
    end
    if (reset) begin // @[DCache.scala 54:26]
      v2_5 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h5 == index_addr) begin // @[DCache.scala 123:26]
      v2_5 <= _d2_T | _GEN_131; // @[DCache.scala 123:26]
    end
    if (reset) begin // @[DCache.scala 54:26]
      v2_6 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h6 == index_addr) begin // @[DCache.scala 123:26]
      v2_6 <= _d2_T | _GEN_131; // @[DCache.scala 123:26]
    end
    if (reset) begin // @[DCache.scala 54:26]
      v2_7 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h7 == index_addr) begin // @[DCache.scala 123:26]
      v2_7 <= _d2_T | _GEN_131; // @[DCache.scala 123:26]
    end
    if (reset) begin // @[DCache.scala 54:26]
      v2_8 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h8 == index_addr) begin // @[DCache.scala 123:26]
      v2_8 <= _d2_T | _GEN_131; // @[DCache.scala 123:26]
    end
    if (reset) begin // @[DCache.scala 54:26]
      v2_9 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h9 == index_addr) begin // @[DCache.scala 123:26]
      v2_9 <= _d2_T | _GEN_131; // @[DCache.scala 123:26]
    end
    if (reset) begin // @[DCache.scala 54:26]
      v2_10 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'ha == index_addr) begin // @[DCache.scala 123:26]
      v2_10 <= _d2_T | _GEN_131; // @[DCache.scala 123:26]
    end
    if (reset) begin // @[DCache.scala 54:26]
      v2_11 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'hb == index_addr) begin // @[DCache.scala 123:26]
      v2_11 <= _d2_T | _GEN_131; // @[DCache.scala 123:26]
    end
    if (reset) begin // @[DCache.scala 54:26]
      v2_12 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'hc == index_addr) begin // @[DCache.scala 123:26]
      v2_12 <= _d2_T | _GEN_131; // @[DCache.scala 123:26]
    end
    if (reset) begin // @[DCache.scala 54:26]
      v2_13 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'hd == index_addr) begin // @[DCache.scala 123:26]
      v2_13 <= _d2_T | _GEN_131; // @[DCache.scala 123:26]
    end
    if (reset) begin // @[DCache.scala 54:26]
      v2_14 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'he == index_addr) begin // @[DCache.scala 123:26]
      v2_14 <= _d2_T | _GEN_131; // @[DCache.scala 123:26]
    end
    if (reset) begin // @[DCache.scala 54:26]
      v2_15 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'hf == index_addr) begin // @[DCache.scala 123:26]
      v2_15 <= _d2_T | _GEN_131; // @[DCache.scala 123:26]
    end
    if (reset) begin // @[DCache.scala 54:26]
      v2_16 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h10 == index_addr) begin // @[DCache.scala 123:26]
      v2_16 <= _d2_T | _GEN_131; // @[DCache.scala 123:26]
    end
    if (reset) begin // @[DCache.scala 54:26]
      v2_17 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h11 == index_addr) begin // @[DCache.scala 123:26]
      v2_17 <= _d2_T | _GEN_131; // @[DCache.scala 123:26]
    end
    if (reset) begin // @[DCache.scala 54:26]
      v2_18 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h12 == index_addr) begin // @[DCache.scala 123:26]
      v2_18 <= _d2_T | _GEN_131; // @[DCache.scala 123:26]
    end
    if (reset) begin // @[DCache.scala 54:26]
      v2_19 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h13 == index_addr) begin // @[DCache.scala 123:26]
      v2_19 <= _d2_T | _GEN_131; // @[DCache.scala 123:26]
    end
    if (reset) begin // @[DCache.scala 54:26]
      v2_20 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h14 == index_addr) begin // @[DCache.scala 123:26]
      v2_20 <= _d2_T | _GEN_131; // @[DCache.scala 123:26]
    end
    if (reset) begin // @[DCache.scala 54:26]
      v2_21 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h15 == index_addr) begin // @[DCache.scala 123:26]
      v2_21 <= _d2_T | _GEN_131; // @[DCache.scala 123:26]
    end
    if (reset) begin // @[DCache.scala 54:26]
      v2_22 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h16 == index_addr) begin // @[DCache.scala 123:26]
      v2_22 <= _d2_T | _GEN_131; // @[DCache.scala 123:26]
    end
    if (reset) begin // @[DCache.scala 54:26]
      v2_23 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h17 == index_addr) begin // @[DCache.scala 123:26]
      v2_23 <= _d2_T | _GEN_131; // @[DCache.scala 123:26]
    end
    if (reset) begin // @[DCache.scala 54:26]
      v2_24 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h18 == index_addr) begin // @[DCache.scala 123:26]
      v2_24 <= _d2_T | _GEN_131; // @[DCache.scala 123:26]
    end
    if (reset) begin // @[DCache.scala 54:26]
      v2_25 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h19 == index_addr) begin // @[DCache.scala 123:26]
      v2_25 <= _d2_T | _GEN_131; // @[DCache.scala 123:26]
    end
    if (reset) begin // @[DCache.scala 54:26]
      v2_26 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h1a == index_addr) begin // @[DCache.scala 123:26]
      v2_26 <= _d2_T | _GEN_131; // @[DCache.scala 123:26]
    end
    if (reset) begin // @[DCache.scala 54:26]
      v2_27 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h1b == index_addr) begin // @[DCache.scala 123:26]
      v2_27 <= _d2_T | _GEN_131; // @[DCache.scala 123:26]
    end
    if (reset) begin // @[DCache.scala 54:26]
      v2_28 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h1c == index_addr) begin // @[DCache.scala 123:26]
      v2_28 <= _d2_T | _GEN_131; // @[DCache.scala 123:26]
    end
    if (reset) begin // @[DCache.scala 54:26]
      v2_29 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h1d == index_addr) begin // @[DCache.scala 123:26]
      v2_29 <= _d2_T | _GEN_131; // @[DCache.scala 123:26]
    end
    if (reset) begin // @[DCache.scala 54:26]
      v2_30 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h1e == index_addr) begin // @[DCache.scala 123:26]
      v2_30 <= _d2_T | _GEN_131; // @[DCache.scala 123:26]
    end
    if (reset) begin // @[DCache.scala 54:26]
      v2_31 <= 1'h0; // @[DCache.scala 54:26]
    end else if (5'h1f == index_addr) begin // @[DCache.scala 123:26]
      v2_31 <= _d2_T | _GEN_131; // @[DCache.scala 123:26]
    end
    if (reset) begin // @[DCache.scala 55:26]
      d2_0 <= 1'h0; // @[DCache.scala 55:26]
    end else if (5'h0 == index_addr) begin // @[DCache.scala 107:20]
      if (update & updateway2) begin // @[DCache.scala 107:26]
        d2_0 <= 1'h0;
      end else begin
        d2_0 <= way2write | _GEN_387;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      d2_1 <= 1'h0; // @[DCache.scala 55:26]
    end else if (5'h1 == index_addr) begin // @[DCache.scala 107:20]
      if (update & updateway2) begin // @[DCache.scala 107:26]
        d2_1 <= 1'h0;
      end else begin
        d2_1 <= way2write | _GEN_387;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      d2_2 <= 1'h0; // @[DCache.scala 55:26]
    end else if (5'h2 == index_addr) begin // @[DCache.scala 107:20]
      if (update & updateway2) begin // @[DCache.scala 107:26]
        d2_2 <= 1'h0;
      end else begin
        d2_2 <= way2write | _GEN_387;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      d2_3 <= 1'h0; // @[DCache.scala 55:26]
    end else if (5'h3 == index_addr) begin // @[DCache.scala 107:20]
      if (update & updateway2) begin // @[DCache.scala 107:26]
        d2_3 <= 1'h0;
      end else begin
        d2_3 <= way2write | _GEN_387;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      d2_4 <= 1'h0; // @[DCache.scala 55:26]
    end else if (5'h4 == index_addr) begin // @[DCache.scala 107:20]
      if (update & updateway2) begin // @[DCache.scala 107:26]
        d2_4 <= 1'h0;
      end else begin
        d2_4 <= way2write | _GEN_387;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      d2_5 <= 1'h0; // @[DCache.scala 55:26]
    end else if (5'h5 == index_addr) begin // @[DCache.scala 107:20]
      if (update & updateway2) begin // @[DCache.scala 107:26]
        d2_5 <= 1'h0;
      end else begin
        d2_5 <= way2write | _GEN_387;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      d2_6 <= 1'h0; // @[DCache.scala 55:26]
    end else if (5'h6 == index_addr) begin // @[DCache.scala 107:20]
      if (update & updateway2) begin // @[DCache.scala 107:26]
        d2_6 <= 1'h0;
      end else begin
        d2_6 <= way2write | _GEN_387;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      d2_7 <= 1'h0; // @[DCache.scala 55:26]
    end else if (5'h7 == index_addr) begin // @[DCache.scala 107:20]
      if (update & updateway2) begin // @[DCache.scala 107:26]
        d2_7 <= 1'h0;
      end else begin
        d2_7 <= way2write | _GEN_387;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      d2_8 <= 1'h0; // @[DCache.scala 55:26]
    end else if (5'h8 == index_addr) begin // @[DCache.scala 107:20]
      if (update & updateway2) begin // @[DCache.scala 107:26]
        d2_8 <= 1'h0;
      end else begin
        d2_8 <= way2write | _GEN_387;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      d2_9 <= 1'h0; // @[DCache.scala 55:26]
    end else if (5'h9 == index_addr) begin // @[DCache.scala 107:20]
      if (update & updateway2) begin // @[DCache.scala 107:26]
        d2_9 <= 1'h0;
      end else begin
        d2_9 <= way2write | _GEN_387;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      d2_10 <= 1'h0; // @[DCache.scala 55:26]
    end else if (5'ha == index_addr) begin // @[DCache.scala 107:20]
      if (update & updateway2) begin // @[DCache.scala 107:26]
        d2_10 <= 1'h0;
      end else begin
        d2_10 <= way2write | _GEN_387;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      d2_11 <= 1'h0; // @[DCache.scala 55:26]
    end else if (5'hb == index_addr) begin // @[DCache.scala 107:20]
      if (update & updateway2) begin // @[DCache.scala 107:26]
        d2_11 <= 1'h0;
      end else begin
        d2_11 <= way2write | _GEN_387;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      d2_12 <= 1'h0; // @[DCache.scala 55:26]
    end else if (5'hc == index_addr) begin // @[DCache.scala 107:20]
      if (update & updateway2) begin // @[DCache.scala 107:26]
        d2_12 <= 1'h0;
      end else begin
        d2_12 <= way2write | _GEN_387;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      d2_13 <= 1'h0; // @[DCache.scala 55:26]
    end else if (5'hd == index_addr) begin // @[DCache.scala 107:20]
      if (update & updateway2) begin // @[DCache.scala 107:26]
        d2_13 <= 1'h0;
      end else begin
        d2_13 <= way2write | _GEN_387;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      d2_14 <= 1'h0; // @[DCache.scala 55:26]
    end else if (5'he == index_addr) begin // @[DCache.scala 107:20]
      if (update & updateway2) begin // @[DCache.scala 107:26]
        d2_14 <= 1'h0;
      end else begin
        d2_14 <= way2write | _GEN_387;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      d2_15 <= 1'h0; // @[DCache.scala 55:26]
    end else if (5'hf == index_addr) begin // @[DCache.scala 107:20]
      if (update & updateway2) begin // @[DCache.scala 107:26]
        d2_15 <= 1'h0;
      end else begin
        d2_15 <= way2write | _GEN_387;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      d2_16 <= 1'h0; // @[DCache.scala 55:26]
    end else if (5'h10 == index_addr) begin // @[DCache.scala 107:20]
      if (update & updateway2) begin // @[DCache.scala 107:26]
        d2_16 <= 1'h0;
      end else begin
        d2_16 <= way2write | _GEN_387;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      d2_17 <= 1'h0; // @[DCache.scala 55:26]
    end else if (5'h11 == index_addr) begin // @[DCache.scala 107:20]
      if (update & updateway2) begin // @[DCache.scala 107:26]
        d2_17 <= 1'h0;
      end else begin
        d2_17 <= way2write | _GEN_387;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      d2_18 <= 1'h0; // @[DCache.scala 55:26]
    end else if (5'h12 == index_addr) begin // @[DCache.scala 107:20]
      if (update & updateway2) begin // @[DCache.scala 107:26]
        d2_18 <= 1'h0;
      end else begin
        d2_18 <= way2write | _GEN_387;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      d2_19 <= 1'h0; // @[DCache.scala 55:26]
    end else if (5'h13 == index_addr) begin // @[DCache.scala 107:20]
      if (update & updateway2) begin // @[DCache.scala 107:26]
        d2_19 <= 1'h0;
      end else begin
        d2_19 <= way2write | _GEN_387;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      d2_20 <= 1'h0; // @[DCache.scala 55:26]
    end else if (5'h14 == index_addr) begin // @[DCache.scala 107:20]
      if (update & updateway2) begin // @[DCache.scala 107:26]
        d2_20 <= 1'h0;
      end else begin
        d2_20 <= way2write | _GEN_387;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      d2_21 <= 1'h0; // @[DCache.scala 55:26]
    end else if (5'h15 == index_addr) begin // @[DCache.scala 107:20]
      if (update & updateway2) begin // @[DCache.scala 107:26]
        d2_21 <= 1'h0;
      end else begin
        d2_21 <= way2write | _GEN_387;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      d2_22 <= 1'h0; // @[DCache.scala 55:26]
    end else if (5'h16 == index_addr) begin // @[DCache.scala 107:20]
      if (update & updateway2) begin // @[DCache.scala 107:26]
        d2_22 <= 1'h0;
      end else begin
        d2_22 <= way2write | _GEN_387;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      d2_23 <= 1'h0; // @[DCache.scala 55:26]
    end else if (5'h17 == index_addr) begin // @[DCache.scala 107:20]
      if (update & updateway2) begin // @[DCache.scala 107:26]
        d2_23 <= 1'h0;
      end else begin
        d2_23 <= way2write | _GEN_387;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      d2_24 <= 1'h0; // @[DCache.scala 55:26]
    end else if (5'h18 == index_addr) begin // @[DCache.scala 107:20]
      if (update & updateway2) begin // @[DCache.scala 107:26]
        d2_24 <= 1'h0;
      end else begin
        d2_24 <= way2write | _GEN_387;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      d2_25 <= 1'h0; // @[DCache.scala 55:26]
    end else if (5'h19 == index_addr) begin // @[DCache.scala 107:20]
      if (update & updateway2) begin // @[DCache.scala 107:26]
        d2_25 <= 1'h0;
      end else begin
        d2_25 <= way2write | _GEN_387;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      d2_26 <= 1'h0; // @[DCache.scala 55:26]
    end else if (5'h1a == index_addr) begin // @[DCache.scala 107:20]
      if (update & updateway2) begin // @[DCache.scala 107:26]
        d2_26 <= 1'h0;
      end else begin
        d2_26 <= way2write | _GEN_387;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      d2_27 <= 1'h0; // @[DCache.scala 55:26]
    end else if (5'h1b == index_addr) begin // @[DCache.scala 107:20]
      if (update & updateway2) begin // @[DCache.scala 107:26]
        d2_27 <= 1'h0;
      end else begin
        d2_27 <= way2write | _GEN_387;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      d2_28 <= 1'h0; // @[DCache.scala 55:26]
    end else if (5'h1c == index_addr) begin // @[DCache.scala 107:20]
      if (update & updateway2) begin // @[DCache.scala 107:26]
        d2_28 <= 1'h0;
      end else begin
        d2_28 <= way2write | _GEN_387;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      d2_29 <= 1'h0; // @[DCache.scala 55:26]
    end else if (5'h1d == index_addr) begin // @[DCache.scala 107:20]
      if (update & updateway2) begin // @[DCache.scala 107:26]
        d2_29 <= 1'h0;
      end else begin
        d2_29 <= way2write | _GEN_387;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      d2_30 <= 1'h0; // @[DCache.scala 55:26]
    end else if (5'h1e == index_addr) begin // @[DCache.scala 107:20]
      if (update & updateway2) begin // @[DCache.scala 107:26]
        d2_30 <= 1'h0;
      end else begin
        d2_30 <= way2write | _GEN_387;
      end
    end
    if (reset) begin // @[DCache.scala 55:26]
      d2_31 <= 1'h0; // @[DCache.scala 55:26]
    end else if (5'h1f == index_addr) begin // @[DCache.scala 107:20]
      if (update & updateway2) begin // @[DCache.scala 107:26]
        d2_31 <= 1'h0;
      end else begin
        d2_31 <= way2write | _GEN_387;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      age2_0 <= 1'h0; // @[DCache.scala 56:26]
    end else if (5'h0 == index_addr) begin // @[DCache.scala 79:22]
      if (_age1_T) begin // @[DCache.scala 79:28]
        age2_0 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 79:28]
        age2_0 <= age2_31; // @[DCache.scala 79:28]
      end else begin
        age2_0 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      age2_1 <= 1'h0; // @[DCache.scala 56:26]
    end else if (5'h1 == index_addr) begin // @[DCache.scala 79:22]
      if (_age1_T) begin // @[DCache.scala 79:28]
        age2_1 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 79:28]
        age2_1 <= age2_31; // @[DCache.scala 79:28]
      end else begin
        age2_1 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      age2_2 <= 1'h0; // @[DCache.scala 56:26]
    end else if (5'h2 == index_addr) begin // @[DCache.scala 79:22]
      if (_age1_T) begin // @[DCache.scala 79:28]
        age2_2 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 79:28]
        age2_2 <= age2_31; // @[DCache.scala 79:28]
      end else begin
        age2_2 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      age2_3 <= 1'h0; // @[DCache.scala 56:26]
    end else if (5'h3 == index_addr) begin // @[DCache.scala 79:22]
      if (_age1_T) begin // @[DCache.scala 79:28]
        age2_3 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 79:28]
        age2_3 <= age2_31; // @[DCache.scala 79:28]
      end else begin
        age2_3 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      age2_4 <= 1'h0; // @[DCache.scala 56:26]
    end else if (5'h4 == index_addr) begin // @[DCache.scala 79:22]
      if (_age1_T) begin // @[DCache.scala 79:28]
        age2_4 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 79:28]
        age2_4 <= age2_31; // @[DCache.scala 79:28]
      end else begin
        age2_4 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      age2_5 <= 1'h0; // @[DCache.scala 56:26]
    end else if (5'h5 == index_addr) begin // @[DCache.scala 79:22]
      if (_age1_T) begin // @[DCache.scala 79:28]
        age2_5 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 79:28]
        age2_5 <= age2_31; // @[DCache.scala 79:28]
      end else begin
        age2_5 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      age2_6 <= 1'h0; // @[DCache.scala 56:26]
    end else if (5'h6 == index_addr) begin // @[DCache.scala 79:22]
      if (_age1_T) begin // @[DCache.scala 79:28]
        age2_6 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 79:28]
        age2_6 <= age2_31; // @[DCache.scala 79:28]
      end else begin
        age2_6 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      age2_7 <= 1'h0; // @[DCache.scala 56:26]
    end else if (5'h7 == index_addr) begin // @[DCache.scala 79:22]
      if (_age1_T) begin // @[DCache.scala 79:28]
        age2_7 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 79:28]
        age2_7 <= age2_31; // @[DCache.scala 79:28]
      end else begin
        age2_7 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      age2_8 <= 1'h0; // @[DCache.scala 56:26]
    end else if (5'h8 == index_addr) begin // @[DCache.scala 79:22]
      if (_age1_T) begin // @[DCache.scala 79:28]
        age2_8 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 79:28]
        age2_8 <= age2_31; // @[DCache.scala 79:28]
      end else begin
        age2_8 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      age2_9 <= 1'h0; // @[DCache.scala 56:26]
    end else if (5'h9 == index_addr) begin // @[DCache.scala 79:22]
      if (_age1_T) begin // @[DCache.scala 79:28]
        age2_9 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 79:28]
        age2_9 <= age2_31; // @[DCache.scala 79:28]
      end else begin
        age2_9 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      age2_10 <= 1'h0; // @[DCache.scala 56:26]
    end else if (5'ha == index_addr) begin // @[DCache.scala 79:22]
      if (_age1_T) begin // @[DCache.scala 79:28]
        age2_10 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 79:28]
        age2_10 <= age2_31; // @[DCache.scala 79:28]
      end else begin
        age2_10 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      age2_11 <= 1'h0; // @[DCache.scala 56:26]
    end else if (5'hb == index_addr) begin // @[DCache.scala 79:22]
      if (_age1_T) begin // @[DCache.scala 79:28]
        age2_11 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 79:28]
        age2_11 <= age2_31; // @[DCache.scala 79:28]
      end else begin
        age2_11 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      age2_12 <= 1'h0; // @[DCache.scala 56:26]
    end else if (5'hc == index_addr) begin // @[DCache.scala 79:22]
      if (_age1_T) begin // @[DCache.scala 79:28]
        age2_12 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 79:28]
        age2_12 <= age2_31; // @[DCache.scala 79:28]
      end else begin
        age2_12 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      age2_13 <= 1'h0; // @[DCache.scala 56:26]
    end else if (5'hd == index_addr) begin // @[DCache.scala 79:22]
      if (_age1_T) begin // @[DCache.scala 79:28]
        age2_13 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 79:28]
        age2_13 <= age2_31; // @[DCache.scala 79:28]
      end else begin
        age2_13 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      age2_14 <= 1'h0; // @[DCache.scala 56:26]
    end else if (5'he == index_addr) begin // @[DCache.scala 79:22]
      if (_age1_T) begin // @[DCache.scala 79:28]
        age2_14 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 79:28]
        age2_14 <= age2_31; // @[DCache.scala 79:28]
      end else begin
        age2_14 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      age2_15 <= 1'h0; // @[DCache.scala 56:26]
    end else if (5'hf == index_addr) begin // @[DCache.scala 79:22]
      if (_age1_T) begin // @[DCache.scala 79:28]
        age2_15 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 79:28]
        age2_15 <= age2_31; // @[DCache.scala 79:28]
      end else begin
        age2_15 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      age2_16 <= 1'h0; // @[DCache.scala 56:26]
    end else if (5'h10 == index_addr) begin // @[DCache.scala 79:22]
      if (_age1_T) begin // @[DCache.scala 79:28]
        age2_16 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 79:28]
        age2_16 <= age2_31; // @[DCache.scala 79:28]
      end else begin
        age2_16 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      age2_17 <= 1'h0; // @[DCache.scala 56:26]
    end else if (5'h11 == index_addr) begin // @[DCache.scala 79:22]
      if (_age1_T) begin // @[DCache.scala 79:28]
        age2_17 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 79:28]
        age2_17 <= age2_31; // @[DCache.scala 79:28]
      end else begin
        age2_17 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      age2_18 <= 1'h0; // @[DCache.scala 56:26]
    end else if (5'h12 == index_addr) begin // @[DCache.scala 79:22]
      if (_age1_T) begin // @[DCache.scala 79:28]
        age2_18 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 79:28]
        age2_18 <= age2_31; // @[DCache.scala 79:28]
      end else begin
        age2_18 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      age2_19 <= 1'h0; // @[DCache.scala 56:26]
    end else if (5'h13 == index_addr) begin // @[DCache.scala 79:22]
      if (_age1_T) begin // @[DCache.scala 79:28]
        age2_19 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 79:28]
        age2_19 <= age2_31; // @[DCache.scala 79:28]
      end else begin
        age2_19 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      age2_20 <= 1'h0; // @[DCache.scala 56:26]
    end else if (5'h14 == index_addr) begin // @[DCache.scala 79:22]
      if (_age1_T) begin // @[DCache.scala 79:28]
        age2_20 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 79:28]
        age2_20 <= age2_31; // @[DCache.scala 79:28]
      end else begin
        age2_20 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      age2_21 <= 1'h0; // @[DCache.scala 56:26]
    end else if (5'h15 == index_addr) begin // @[DCache.scala 79:22]
      if (_age1_T) begin // @[DCache.scala 79:28]
        age2_21 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 79:28]
        age2_21 <= age2_31; // @[DCache.scala 79:28]
      end else begin
        age2_21 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      age2_22 <= 1'h0; // @[DCache.scala 56:26]
    end else if (5'h16 == index_addr) begin // @[DCache.scala 79:22]
      if (_age1_T) begin // @[DCache.scala 79:28]
        age2_22 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 79:28]
        age2_22 <= age2_31; // @[DCache.scala 79:28]
      end else begin
        age2_22 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      age2_23 <= 1'h0; // @[DCache.scala 56:26]
    end else if (5'h17 == index_addr) begin // @[DCache.scala 79:22]
      if (_age1_T) begin // @[DCache.scala 79:28]
        age2_23 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 79:28]
        age2_23 <= age2_31; // @[DCache.scala 79:28]
      end else begin
        age2_23 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      age2_24 <= 1'h0; // @[DCache.scala 56:26]
    end else if (5'h18 == index_addr) begin // @[DCache.scala 79:22]
      if (_age1_T) begin // @[DCache.scala 79:28]
        age2_24 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 79:28]
        age2_24 <= age2_31; // @[DCache.scala 79:28]
      end else begin
        age2_24 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      age2_25 <= 1'h0; // @[DCache.scala 56:26]
    end else if (5'h19 == index_addr) begin // @[DCache.scala 79:22]
      if (_age1_T) begin // @[DCache.scala 79:28]
        age2_25 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 79:28]
        age2_25 <= age2_31; // @[DCache.scala 79:28]
      end else begin
        age2_25 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      age2_26 <= 1'h0; // @[DCache.scala 56:26]
    end else if (5'h1a == index_addr) begin // @[DCache.scala 79:22]
      if (_age1_T) begin // @[DCache.scala 79:28]
        age2_26 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 79:28]
        age2_26 <= age2_31; // @[DCache.scala 79:28]
      end else begin
        age2_26 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      age2_27 <= 1'h0; // @[DCache.scala 56:26]
    end else if (5'h1b == index_addr) begin // @[DCache.scala 79:22]
      if (_age1_T) begin // @[DCache.scala 79:28]
        age2_27 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 79:28]
        age2_27 <= age2_31; // @[DCache.scala 79:28]
      end else begin
        age2_27 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      age2_28 <= 1'h0; // @[DCache.scala 56:26]
    end else if (5'h1c == index_addr) begin // @[DCache.scala 79:22]
      if (_age1_T) begin // @[DCache.scala 79:28]
        age2_28 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 79:28]
        age2_28 <= age2_31; // @[DCache.scala 79:28]
      end else begin
        age2_28 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      age2_29 <= 1'h0; // @[DCache.scala 56:26]
    end else if (5'h1d == index_addr) begin // @[DCache.scala 79:22]
      if (_age1_T) begin // @[DCache.scala 79:28]
        age2_29 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 79:28]
        age2_29 <= age2_31; // @[DCache.scala 79:28]
      end else begin
        age2_29 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      age2_30 <= 1'h0; // @[DCache.scala 56:26]
    end else if (5'h1e == index_addr) begin // @[DCache.scala 79:22]
      if (_age1_T) begin // @[DCache.scala 79:28]
        age2_30 <= hit2;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 79:28]
        age2_30 <= age2_31; // @[DCache.scala 79:28]
      end else begin
        age2_30 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 56:26]
      age2_31 <= 1'h0; // @[DCache.scala 56:26]
    end else if (5'h1f == index_addr) begin // @[DCache.scala 79:22]
      if (_age1_T) begin // @[DCache.scala 79:28]
        age2_31 <= hit2;
      end else if (!(5'h1f == index_addr)) begin // @[DCache.scala 79:28]
        age2_31 <= _GEN_290;
      end
    end
    if (reset) begin // @[DCache.scala 57:26]
      tag2_0 <= 53'h0; // @[DCache.scala 57:26]
    end else if (5'h0 == index_addr) begin // @[DCache.scala 122:26]
      if (_d2_T) begin // @[DCache.scala 122:32]
        tag2_0 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 61:28]
        tag2_0 <= tag2_31; // @[DCache.scala 61:28]
      end else begin
        tag2_0 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 57:26]
      tag2_1 <= 53'h0; // @[DCache.scala 57:26]
    end else if (5'h1 == index_addr) begin // @[DCache.scala 122:26]
      if (_d2_T) begin // @[DCache.scala 122:32]
        tag2_1 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 61:28]
        tag2_1 <= tag2_31; // @[DCache.scala 61:28]
      end else begin
        tag2_1 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 57:26]
      tag2_2 <= 53'h0; // @[DCache.scala 57:26]
    end else if (5'h2 == index_addr) begin // @[DCache.scala 122:26]
      if (_d2_T) begin // @[DCache.scala 122:32]
        tag2_2 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 61:28]
        tag2_2 <= tag2_31; // @[DCache.scala 61:28]
      end else begin
        tag2_2 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 57:26]
      tag2_3 <= 53'h0; // @[DCache.scala 57:26]
    end else if (5'h3 == index_addr) begin // @[DCache.scala 122:26]
      if (_d2_T) begin // @[DCache.scala 122:32]
        tag2_3 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 61:28]
        tag2_3 <= tag2_31; // @[DCache.scala 61:28]
      end else begin
        tag2_3 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 57:26]
      tag2_4 <= 53'h0; // @[DCache.scala 57:26]
    end else if (5'h4 == index_addr) begin // @[DCache.scala 122:26]
      if (_d2_T) begin // @[DCache.scala 122:32]
        tag2_4 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 61:28]
        tag2_4 <= tag2_31; // @[DCache.scala 61:28]
      end else begin
        tag2_4 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 57:26]
      tag2_5 <= 53'h0; // @[DCache.scala 57:26]
    end else if (5'h5 == index_addr) begin // @[DCache.scala 122:26]
      if (_d2_T) begin // @[DCache.scala 122:32]
        tag2_5 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 61:28]
        tag2_5 <= tag2_31; // @[DCache.scala 61:28]
      end else begin
        tag2_5 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 57:26]
      tag2_6 <= 53'h0; // @[DCache.scala 57:26]
    end else if (5'h6 == index_addr) begin // @[DCache.scala 122:26]
      if (_d2_T) begin // @[DCache.scala 122:32]
        tag2_6 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 61:28]
        tag2_6 <= tag2_31; // @[DCache.scala 61:28]
      end else begin
        tag2_6 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 57:26]
      tag2_7 <= 53'h0; // @[DCache.scala 57:26]
    end else if (5'h7 == index_addr) begin // @[DCache.scala 122:26]
      if (_d2_T) begin // @[DCache.scala 122:32]
        tag2_7 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 61:28]
        tag2_7 <= tag2_31; // @[DCache.scala 61:28]
      end else begin
        tag2_7 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 57:26]
      tag2_8 <= 53'h0; // @[DCache.scala 57:26]
    end else if (5'h8 == index_addr) begin // @[DCache.scala 122:26]
      if (_d2_T) begin // @[DCache.scala 122:32]
        tag2_8 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 61:28]
        tag2_8 <= tag2_31; // @[DCache.scala 61:28]
      end else begin
        tag2_8 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 57:26]
      tag2_9 <= 53'h0; // @[DCache.scala 57:26]
    end else if (5'h9 == index_addr) begin // @[DCache.scala 122:26]
      if (_d2_T) begin // @[DCache.scala 122:32]
        tag2_9 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 61:28]
        tag2_9 <= tag2_31; // @[DCache.scala 61:28]
      end else begin
        tag2_9 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 57:26]
      tag2_10 <= 53'h0; // @[DCache.scala 57:26]
    end else if (5'ha == index_addr) begin // @[DCache.scala 122:26]
      if (_d2_T) begin // @[DCache.scala 122:32]
        tag2_10 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 61:28]
        tag2_10 <= tag2_31; // @[DCache.scala 61:28]
      end else begin
        tag2_10 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 57:26]
      tag2_11 <= 53'h0; // @[DCache.scala 57:26]
    end else if (5'hb == index_addr) begin // @[DCache.scala 122:26]
      if (_d2_T) begin // @[DCache.scala 122:32]
        tag2_11 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 61:28]
        tag2_11 <= tag2_31; // @[DCache.scala 61:28]
      end else begin
        tag2_11 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 57:26]
      tag2_12 <= 53'h0; // @[DCache.scala 57:26]
    end else if (5'hc == index_addr) begin // @[DCache.scala 122:26]
      if (_d2_T) begin // @[DCache.scala 122:32]
        tag2_12 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 61:28]
        tag2_12 <= tag2_31; // @[DCache.scala 61:28]
      end else begin
        tag2_12 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 57:26]
      tag2_13 <= 53'h0; // @[DCache.scala 57:26]
    end else if (5'hd == index_addr) begin // @[DCache.scala 122:26]
      if (_d2_T) begin // @[DCache.scala 122:32]
        tag2_13 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 61:28]
        tag2_13 <= tag2_31; // @[DCache.scala 61:28]
      end else begin
        tag2_13 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 57:26]
      tag2_14 <= 53'h0; // @[DCache.scala 57:26]
    end else if (5'he == index_addr) begin // @[DCache.scala 122:26]
      if (_d2_T) begin // @[DCache.scala 122:32]
        tag2_14 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 61:28]
        tag2_14 <= tag2_31; // @[DCache.scala 61:28]
      end else begin
        tag2_14 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 57:26]
      tag2_15 <= 53'h0; // @[DCache.scala 57:26]
    end else if (5'hf == index_addr) begin // @[DCache.scala 122:26]
      if (_d2_T) begin // @[DCache.scala 122:32]
        tag2_15 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 61:28]
        tag2_15 <= tag2_31; // @[DCache.scala 61:28]
      end else begin
        tag2_15 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 57:26]
      tag2_16 <= 53'h0; // @[DCache.scala 57:26]
    end else if (5'h10 == index_addr) begin // @[DCache.scala 122:26]
      if (_d2_T) begin // @[DCache.scala 122:32]
        tag2_16 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 61:28]
        tag2_16 <= tag2_31; // @[DCache.scala 61:28]
      end else begin
        tag2_16 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 57:26]
      tag2_17 <= 53'h0; // @[DCache.scala 57:26]
    end else if (5'h11 == index_addr) begin // @[DCache.scala 122:26]
      if (_d2_T) begin // @[DCache.scala 122:32]
        tag2_17 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 61:28]
        tag2_17 <= tag2_31; // @[DCache.scala 61:28]
      end else begin
        tag2_17 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 57:26]
      tag2_18 <= 53'h0; // @[DCache.scala 57:26]
    end else if (5'h12 == index_addr) begin // @[DCache.scala 122:26]
      if (_d2_T) begin // @[DCache.scala 122:32]
        tag2_18 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 61:28]
        tag2_18 <= tag2_31; // @[DCache.scala 61:28]
      end else begin
        tag2_18 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 57:26]
      tag2_19 <= 53'h0; // @[DCache.scala 57:26]
    end else if (5'h13 == index_addr) begin // @[DCache.scala 122:26]
      if (_d2_T) begin // @[DCache.scala 122:32]
        tag2_19 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 61:28]
        tag2_19 <= tag2_31; // @[DCache.scala 61:28]
      end else begin
        tag2_19 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 57:26]
      tag2_20 <= 53'h0; // @[DCache.scala 57:26]
    end else if (5'h14 == index_addr) begin // @[DCache.scala 122:26]
      if (_d2_T) begin // @[DCache.scala 122:32]
        tag2_20 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 61:28]
        tag2_20 <= tag2_31; // @[DCache.scala 61:28]
      end else begin
        tag2_20 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 57:26]
      tag2_21 <= 53'h0; // @[DCache.scala 57:26]
    end else if (5'h15 == index_addr) begin // @[DCache.scala 122:26]
      if (_d2_T) begin // @[DCache.scala 122:32]
        tag2_21 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 61:28]
        tag2_21 <= tag2_31; // @[DCache.scala 61:28]
      end else begin
        tag2_21 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 57:26]
      tag2_22 <= 53'h0; // @[DCache.scala 57:26]
    end else if (5'h16 == index_addr) begin // @[DCache.scala 122:26]
      if (_d2_T) begin // @[DCache.scala 122:32]
        tag2_22 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 61:28]
        tag2_22 <= tag2_31; // @[DCache.scala 61:28]
      end else begin
        tag2_22 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 57:26]
      tag2_23 <= 53'h0; // @[DCache.scala 57:26]
    end else if (5'h17 == index_addr) begin // @[DCache.scala 122:26]
      if (_d2_T) begin // @[DCache.scala 122:32]
        tag2_23 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 61:28]
        tag2_23 <= tag2_31; // @[DCache.scala 61:28]
      end else begin
        tag2_23 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 57:26]
      tag2_24 <= 53'h0; // @[DCache.scala 57:26]
    end else if (5'h18 == index_addr) begin // @[DCache.scala 122:26]
      if (_d2_T) begin // @[DCache.scala 122:32]
        tag2_24 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 61:28]
        tag2_24 <= tag2_31; // @[DCache.scala 61:28]
      end else begin
        tag2_24 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 57:26]
      tag2_25 <= 53'h0; // @[DCache.scala 57:26]
    end else if (5'h19 == index_addr) begin // @[DCache.scala 122:26]
      if (_d2_T) begin // @[DCache.scala 122:32]
        tag2_25 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 61:28]
        tag2_25 <= tag2_31; // @[DCache.scala 61:28]
      end else begin
        tag2_25 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 57:26]
      tag2_26 <= 53'h0; // @[DCache.scala 57:26]
    end else if (5'h1a == index_addr) begin // @[DCache.scala 122:26]
      if (_d2_T) begin // @[DCache.scala 122:32]
        tag2_26 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 61:28]
        tag2_26 <= tag2_31; // @[DCache.scala 61:28]
      end else begin
        tag2_26 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 57:26]
      tag2_27 <= 53'h0; // @[DCache.scala 57:26]
    end else if (5'h1b == index_addr) begin // @[DCache.scala 122:26]
      if (_d2_T) begin // @[DCache.scala 122:32]
        tag2_27 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 61:28]
        tag2_27 <= tag2_31; // @[DCache.scala 61:28]
      end else begin
        tag2_27 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 57:26]
      tag2_28 <= 53'h0; // @[DCache.scala 57:26]
    end else if (5'h1c == index_addr) begin // @[DCache.scala 122:26]
      if (_d2_T) begin // @[DCache.scala 122:32]
        tag2_28 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 61:28]
        tag2_28 <= tag2_31; // @[DCache.scala 61:28]
      end else begin
        tag2_28 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 57:26]
      tag2_29 <= 53'h0; // @[DCache.scala 57:26]
    end else if (5'h1d == index_addr) begin // @[DCache.scala 122:26]
      if (_d2_T) begin // @[DCache.scala 122:32]
        tag2_29 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 61:28]
        tag2_29 <= tag2_31; // @[DCache.scala 61:28]
      end else begin
        tag2_29 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 57:26]
      tag2_30 <= 53'h0; // @[DCache.scala 57:26]
    end else if (5'h1e == index_addr) begin // @[DCache.scala 122:26]
      if (_d2_T) begin // @[DCache.scala 122:32]
        tag2_30 <= tag_addr;
      end else if (5'h1f == index_addr) begin // @[DCache.scala 61:28]
        tag2_30 <= tag2_31; // @[DCache.scala 61:28]
      end else begin
        tag2_30 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 57:26]
      tag2_31 <= 53'h0; // @[DCache.scala 57:26]
    end else if (5'h1f == index_addr) begin // @[DCache.scala 122:26]
      if (_d2_T) begin // @[DCache.scala 122:32]
        tag2_31 <= tag_addr;
      end else if (!(5'h1f == index_addr)) begin // @[DCache.scala 61:28]
        tag2_31 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCache.scala 58:26]
      block2_0 <= 512'h0; // @[DCache.scala 58:26]
    end else if (5'h0 == index_addr) begin // @[DCache.scala 121:26]
      if (_d2_T) begin // @[DCache.scala 121:32]
        block2_0 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 121:72]
        block2_0 <= block2_after_write;
      end else begin
        block2_0 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 58:26]
      block2_1 <= 512'h0; // @[DCache.scala 58:26]
    end else if (5'h1 == index_addr) begin // @[DCache.scala 121:26]
      if (_d2_T) begin // @[DCache.scala 121:32]
        block2_1 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 121:72]
        block2_1 <= block2_after_write;
      end else begin
        block2_1 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 58:26]
      block2_2 <= 512'h0; // @[DCache.scala 58:26]
    end else if (5'h2 == index_addr) begin // @[DCache.scala 121:26]
      if (_d2_T) begin // @[DCache.scala 121:32]
        block2_2 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 121:72]
        block2_2 <= block2_after_write;
      end else begin
        block2_2 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 58:26]
      block2_3 <= 512'h0; // @[DCache.scala 58:26]
    end else if (5'h3 == index_addr) begin // @[DCache.scala 121:26]
      if (_d2_T) begin // @[DCache.scala 121:32]
        block2_3 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 121:72]
        block2_3 <= block2_after_write;
      end else begin
        block2_3 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 58:26]
      block2_4 <= 512'h0; // @[DCache.scala 58:26]
    end else if (5'h4 == index_addr) begin // @[DCache.scala 121:26]
      if (_d2_T) begin // @[DCache.scala 121:32]
        block2_4 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 121:72]
        block2_4 <= block2_after_write;
      end else begin
        block2_4 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 58:26]
      block2_5 <= 512'h0; // @[DCache.scala 58:26]
    end else if (5'h5 == index_addr) begin // @[DCache.scala 121:26]
      if (_d2_T) begin // @[DCache.scala 121:32]
        block2_5 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 121:72]
        block2_5 <= block2_after_write;
      end else begin
        block2_5 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 58:26]
      block2_6 <= 512'h0; // @[DCache.scala 58:26]
    end else if (5'h6 == index_addr) begin // @[DCache.scala 121:26]
      if (_d2_T) begin // @[DCache.scala 121:32]
        block2_6 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 121:72]
        block2_6 <= block2_after_write;
      end else begin
        block2_6 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 58:26]
      block2_7 <= 512'h0; // @[DCache.scala 58:26]
    end else if (5'h7 == index_addr) begin // @[DCache.scala 121:26]
      if (_d2_T) begin // @[DCache.scala 121:32]
        block2_7 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 121:72]
        block2_7 <= block2_after_write;
      end else begin
        block2_7 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 58:26]
      block2_8 <= 512'h0; // @[DCache.scala 58:26]
    end else if (5'h8 == index_addr) begin // @[DCache.scala 121:26]
      if (_d2_T) begin // @[DCache.scala 121:32]
        block2_8 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 121:72]
        block2_8 <= block2_after_write;
      end else begin
        block2_8 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 58:26]
      block2_9 <= 512'h0; // @[DCache.scala 58:26]
    end else if (5'h9 == index_addr) begin // @[DCache.scala 121:26]
      if (_d2_T) begin // @[DCache.scala 121:32]
        block2_9 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 121:72]
        block2_9 <= block2_after_write;
      end else begin
        block2_9 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 58:26]
      block2_10 <= 512'h0; // @[DCache.scala 58:26]
    end else if (5'ha == index_addr) begin // @[DCache.scala 121:26]
      if (_d2_T) begin // @[DCache.scala 121:32]
        block2_10 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 121:72]
        block2_10 <= block2_after_write;
      end else begin
        block2_10 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 58:26]
      block2_11 <= 512'h0; // @[DCache.scala 58:26]
    end else if (5'hb == index_addr) begin // @[DCache.scala 121:26]
      if (_d2_T) begin // @[DCache.scala 121:32]
        block2_11 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 121:72]
        block2_11 <= block2_after_write;
      end else begin
        block2_11 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 58:26]
      block2_12 <= 512'h0; // @[DCache.scala 58:26]
    end else if (5'hc == index_addr) begin // @[DCache.scala 121:26]
      if (_d2_T) begin // @[DCache.scala 121:32]
        block2_12 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 121:72]
        block2_12 <= block2_after_write;
      end else begin
        block2_12 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 58:26]
      block2_13 <= 512'h0; // @[DCache.scala 58:26]
    end else if (5'hd == index_addr) begin // @[DCache.scala 121:26]
      if (_d2_T) begin // @[DCache.scala 121:32]
        block2_13 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 121:72]
        block2_13 <= block2_after_write;
      end else begin
        block2_13 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 58:26]
      block2_14 <= 512'h0; // @[DCache.scala 58:26]
    end else if (5'he == index_addr) begin // @[DCache.scala 121:26]
      if (_d2_T) begin // @[DCache.scala 121:32]
        block2_14 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 121:72]
        block2_14 <= block2_after_write;
      end else begin
        block2_14 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 58:26]
      block2_15 <= 512'h0; // @[DCache.scala 58:26]
    end else if (5'hf == index_addr) begin // @[DCache.scala 121:26]
      if (_d2_T) begin // @[DCache.scala 121:32]
        block2_15 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 121:72]
        block2_15 <= block2_after_write;
      end else begin
        block2_15 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 58:26]
      block2_16 <= 512'h0; // @[DCache.scala 58:26]
    end else if (5'h10 == index_addr) begin // @[DCache.scala 121:26]
      if (_d2_T) begin // @[DCache.scala 121:32]
        block2_16 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 121:72]
        block2_16 <= block2_after_write;
      end else begin
        block2_16 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 58:26]
      block2_17 <= 512'h0; // @[DCache.scala 58:26]
    end else if (5'h11 == index_addr) begin // @[DCache.scala 121:26]
      if (_d2_T) begin // @[DCache.scala 121:32]
        block2_17 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 121:72]
        block2_17 <= block2_after_write;
      end else begin
        block2_17 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 58:26]
      block2_18 <= 512'h0; // @[DCache.scala 58:26]
    end else if (5'h12 == index_addr) begin // @[DCache.scala 121:26]
      if (_d2_T) begin // @[DCache.scala 121:32]
        block2_18 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 121:72]
        block2_18 <= block2_after_write;
      end else begin
        block2_18 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 58:26]
      block2_19 <= 512'h0; // @[DCache.scala 58:26]
    end else if (5'h13 == index_addr) begin // @[DCache.scala 121:26]
      if (_d2_T) begin // @[DCache.scala 121:32]
        block2_19 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 121:72]
        block2_19 <= block2_after_write;
      end else begin
        block2_19 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 58:26]
      block2_20 <= 512'h0; // @[DCache.scala 58:26]
    end else if (5'h14 == index_addr) begin // @[DCache.scala 121:26]
      if (_d2_T) begin // @[DCache.scala 121:32]
        block2_20 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 121:72]
        block2_20 <= block2_after_write;
      end else begin
        block2_20 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 58:26]
      block2_21 <= 512'h0; // @[DCache.scala 58:26]
    end else if (5'h15 == index_addr) begin // @[DCache.scala 121:26]
      if (_d2_T) begin // @[DCache.scala 121:32]
        block2_21 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 121:72]
        block2_21 <= block2_after_write;
      end else begin
        block2_21 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 58:26]
      block2_22 <= 512'h0; // @[DCache.scala 58:26]
    end else if (5'h16 == index_addr) begin // @[DCache.scala 121:26]
      if (_d2_T) begin // @[DCache.scala 121:32]
        block2_22 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 121:72]
        block2_22 <= block2_after_write;
      end else begin
        block2_22 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 58:26]
      block2_23 <= 512'h0; // @[DCache.scala 58:26]
    end else if (5'h17 == index_addr) begin // @[DCache.scala 121:26]
      if (_d2_T) begin // @[DCache.scala 121:32]
        block2_23 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 121:72]
        block2_23 <= block2_after_write;
      end else begin
        block2_23 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 58:26]
      block2_24 <= 512'h0; // @[DCache.scala 58:26]
    end else if (5'h18 == index_addr) begin // @[DCache.scala 121:26]
      if (_d2_T) begin // @[DCache.scala 121:32]
        block2_24 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 121:72]
        block2_24 <= block2_after_write;
      end else begin
        block2_24 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 58:26]
      block2_25 <= 512'h0; // @[DCache.scala 58:26]
    end else if (5'h19 == index_addr) begin // @[DCache.scala 121:26]
      if (_d2_T) begin // @[DCache.scala 121:32]
        block2_25 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 121:72]
        block2_25 <= block2_after_write;
      end else begin
        block2_25 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 58:26]
      block2_26 <= 512'h0; // @[DCache.scala 58:26]
    end else if (5'h1a == index_addr) begin // @[DCache.scala 121:26]
      if (_d2_T) begin // @[DCache.scala 121:32]
        block2_26 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 121:72]
        block2_26 <= block2_after_write;
      end else begin
        block2_26 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 58:26]
      block2_27 <= 512'h0; // @[DCache.scala 58:26]
    end else if (5'h1b == index_addr) begin // @[DCache.scala 121:26]
      if (_d2_T) begin // @[DCache.scala 121:32]
        block2_27 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 121:72]
        block2_27 <= block2_after_write;
      end else begin
        block2_27 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 58:26]
      block2_28 <= 512'h0; // @[DCache.scala 58:26]
    end else if (5'h1c == index_addr) begin // @[DCache.scala 121:26]
      if (_d2_T) begin // @[DCache.scala 121:32]
        block2_28 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 121:72]
        block2_28 <= block2_after_write;
      end else begin
        block2_28 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 58:26]
      block2_29 <= 512'h0; // @[DCache.scala 58:26]
    end else if (5'h1d == index_addr) begin // @[DCache.scala 121:26]
      if (_d2_T) begin // @[DCache.scala 121:32]
        block2_29 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 121:72]
        block2_29 <= block2_after_write;
      end else begin
        block2_29 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 58:26]
      block2_30 <= 512'h0; // @[DCache.scala 58:26]
    end else if (5'h1e == index_addr) begin // @[DCache.scala 121:26]
      if (_d2_T) begin // @[DCache.scala 121:32]
        block2_30 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 121:72]
        block2_30 <= block2_after_write;
      end else begin
        block2_30 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 58:26]
      block2_31 <= 512'h0; // @[DCache.scala 58:26]
    end else if (5'h1f == index_addr) begin // @[DCache.scala 121:26]
      if (_d2_T) begin // @[DCache.scala 121:32]
        block2_31 <= io_axi_rdata;
      end else if (way2write) begin // @[DCache.scala 121:72]
        block2_31 <= block2_after_write;
      end else begin
        block2_31 <= _GEN_195;
      end
    end
    if (reset) begin // @[DCache.scala 66:24]
      state <= 2'h0; // @[DCache.scala 66:24]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (miss & ~not_en_yet) begin // @[DCache.scala 90:39]
        if (dirty) begin // @[DCache.scala 90:52]
          state <= 2'h1;
        end else begin
          state <= 2'h2;
        end
      end
    end else if (_T_3) begin // @[Conditional.scala 39:67]
      if (io_axi_wdone) begin // @[DCache.scala 94:32]
        state <= 2'h2; // @[DCache.scala 94:39]
      end
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      state <= _GEN_390;
    end
    not_en_yet <= reset | _not_en_yet_T; // @[DCache.scala 71:30 DCache.scala 71:30 DCache.scala 72:21]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  op = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  addr = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  wdata = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  wm = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  v1_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  v1_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  v1_2 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  v1_3 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  v1_4 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  v1_5 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  v1_6 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  v1_7 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  v1_8 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  v1_9 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  v1_10 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  v1_11 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  v1_12 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  v1_13 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  v1_14 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  v1_15 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  v1_16 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  v1_17 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  v1_18 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  v1_19 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  v1_20 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  v1_21 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  v1_22 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  v1_23 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  v1_24 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  v1_25 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  v1_26 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  v1_27 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  v1_28 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  v1_29 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  v1_30 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  v1_31 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  d1_0 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  d1_1 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  d1_2 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  d1_3 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  d1_4 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  d1_5 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  d1_6 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  d1_7 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  d1_8 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  d1_9 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  d1_10 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  d1_11 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  d1_12 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  d1_13 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  d1_14 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  d1_15 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  d1_16 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  d1_17 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  d1_18 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  d1_19 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  d1_20 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  d1_21 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  d1_22 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  d1_23 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  d1_24 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  d1_25 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  d1_26 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  d1_27 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  d1_28 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  d1_29 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  d1_30 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  d1_31 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  age1_0 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  age1_1 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  age1_2 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  age1_3 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  age1_4 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  age1_5 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  age1_6 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  age1_7 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  age1_8 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  age1_9 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  age1_10 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  age1_11 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  age1_12 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  age1_13 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  age1_14 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  age1_15 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  age1_16 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  age1_17 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  age1_18 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  age1_19 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  age1_20 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  age1_21 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  age1_22 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  age1_23 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  age1_24 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  age1_25 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  age1_26 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  age1_27 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  age1_28 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  age1_29 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  age1_30 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  age1_31 = _RAND_99[0:0];
  _RAND_100 = {2{`RANDOM}};
  tag1_0 = _RAND_100[52:0];
  _RAND_101 = {2{`RANDOM}};
  tag1_1 = _RAND_101[52:0];
  _RAND_102 = {2{`RANDOM}};
  tag1_2 = _RAND_102[52:0];
  _RAND_103 = {2{`RANDOM}};
  tag1_3 = _RAND_103[52:0];
  _RAND_104 = {2{`RANDOM}};
  tag1_4 = _RAND_104[52:0];
  _RAND_105 = {2{`RANDOM}};
  tag1_5 = _RAND_105[52:0];
  _RAND_106 = {2{`RANDOM}};
  tag1_6 = _RAND_106[52:0];
  _RAND_107 = {2{`RANDOM}};
  tag1_7 = _RAND_107[52:0];
  _RAND_108 = {2{`RANDOM}};
  tag1_8 = _RAND_108[52:0];
  _RAND_109 = {2{`RANDOM}};
  tag1_9 = _RAND_109[52:0];
  _RAND_110 = {2{`RANDOM}};
  tag1_10 = _RAND_110[52:0];
  _RAND_111 = {2{`RANDOM}};
  tag1_11 = _RAND_111[52:0];
  _RAND_112 = {2{`RANDOM}};
  tag1_12 = _RAND_112[52:0];
  _RAND_113 = {2{`RANDOM}};
  tag1_13 = _RAND_113[52:0];
  _RAND_114 = {2{`RANDOM}};
  tag1_14 = _RAND_114[52:0];
  _RAND_115 = {2{`RANDOM}};
  tag1_15 = _RAND_115[52:0];
  _RAND_116 = {2{`RANDOM}};
  tag1_16 = _RAND_116[52:0];
  _RAND_117 = {2{`RANDOM}};
  tag1_17 = _RAND_117[52:0];
  _RAND_118 = {2{`RANDOM}};
  tag1_18 = _RAND_118[52:0];
  _RAND_119 = {2{`RANDOM}};
  tag1_19 = _RAND_119[52:0];
  _RAND_120 = {2{`RANDOM}};
  tag1_20 = _RAND_120[52:0];
  _RAND_121 = {2{`RANDOM}};
  tag1_21 = _RAND_121[52:0];
  _RAND_122 = {2{`RANDOM}};
  tag1_22 = _RAND_122[52:0];
  _RAND_123 = {2{`RANDOM}};
  tag1_23 = _RAND_123[52:0];
  _RAND_124 = {2{`RANDOM}};
  tag1_24 = _RAND_124[52:0];
  _RAND_125 = {2{`RANDOM}};
  tag1_25 = _RAND_125[52:0];
  _RAND_126 = {2{`RANDOM}};
  tag1_26 = _RAND_126[52:0];
  _RAND_127 = {2{`RANDOM}};
  tag1_27 = _RAND_127[52:0];
  _RAND_128 = {2{`RANDOM}};
  tag1_28 = _RAND_128[52:0];
  _RAND_129 = {2{`RANDOM}};
  tag1_29 = _RAND_129[52:0];
  _RAND_130 = {2{`RANDOM}};
  tag1_30 = _RAND_130[52:0];
  _RAND_131 = {2{`RANDOM}};
  tag1_31 = _RAND_131[52:0];
  _RAND_132 = {16{`RANDOM}};
  block1_0 = _RAND_132[511:0];
  _RAND_133 = {16{`RANDOM}};
  block1_1 = _RAND_133[511:0];
  _RAND_134 = {16{`RANDOM}};
  block1_2 = _RAND_134[511:0];
  _RAND_135 = {16{`RANDOM}};
  block1_3 = _RAND_135[511:0];
  _RAND_136 = {16{`RANDOM}};
  block1_4 = _RAND_136[511:0];
  _RAND_137 = {16{`RANDOM}};
  block1_5 = _RAND_137[511:0];
  _RAND_138 = {16{`RANDOM}};
  block1_6 = _RAND_138[511:0];
  _RAND_139 = {16{`RANDOM}};
  block1_7 = _RAND_139[511:0];
  _RAND_140 = {16{`RANDOM}};
  block1_8 = _RAND_140[511:0];
  _RAND_141 = {16{`RANDOM}};
  block1_9 = _RAND_141[511:0];
  _RAND_142 = {16{`RANDOM}};
  block1_10 = _RAND_142[511:0];
  _RAND_143 = {16{`RANDOM}};
  block1_11 = _RAND_143[511:0];
  _RAND_144 = {16{`RANDOM}};
  block1_12 = _RAND_144[511:0];
  _RAND_145 = {16{`RANDOM}};
  block1_13 = _RAND_145[511:0];
  _RAND_146 = {16{`RANDOM}};
  block1_14 = _RAND_146[511:0];
  _RAND_147 = {16{`RANDOM}};
  block1_15 = _RAND_147[511:0];
  _RAND_148 = {16{`RANDOM}};
  block1_16 = _RAND_148[511:0];
  _RAND_149 = {16{`RANDOM}};
  block1_17 = _RAND_149[511:0];
  _RAND_150 = {16{`RANDOM}};
  block1_18 = _RAND_150[511:0];
  _RAND_151 = {16{`RANDOM}};
  block1_19 = _RAND_151[511:0];
  _RAND_152 = {16{`RANDOM}};
  block1_20 = _RAND_152[511:0];
  _RAND_153 = {16{`RANDOM}};
  block1_21 = _RAND_153[511:0];
  _RAND_154 = {16{`RANDOM}};
  block1_22 = _RAND_154[511:0];
  _RAND_155 = {16{`RANDOM}};
  block1_23 = _RAND_155[511:0];
  _RAND_156 = {16{`RANDOM}};
  block1_24 = _RAND_156[511:0];
  _RAND_157 = {16{`RANDOM}};
  block1_25 = _RAND_157[511:0];
  _RAND_158 = {16{`RANDOM}};
  block1_26 = _RAND_158[511:0];
  _RAND_159 = {16{`RANDOM}};
  block1_27 = _RAND_159[511:0];
  _RAND_160 = {16{`RANDOM}};
  block1_28 = _RAND_160[511:0];
  _RAND_161 = {16{`RANDOM}};
  block1_29 = _RAND_161[511:0];
  _RAND_162 = {16{`RANDOM}};
  block1_30 = _RAND_162[511:0];
  _RAND_163 = {16{`RANDOM}};
  block1_31 = _RAND_163[511:0];
  _RAND_164 = {1{`RANDOM}};
  v2_0 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  v2_1 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  v2_2 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  v2_3 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  v2_4 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  v2_5 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  v2_6 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  v2_7 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  v2_8 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  v2_9 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  v2_10 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  v2_11 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  v2_12 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  v2_13 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  v2_14 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  v2_15 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  v2_16 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  v2_17 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  v2_18 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  v2_19 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  v2_20 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  v2_21 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  v2_22 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  v2_23 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  v2_24 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  v2_25 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  v2_26 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  v2_27 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  v2_28 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  v2_29 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  v2_30 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  v2_31 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  d2_0 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  d2_1 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  d2_2 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  d2_3 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  d2_4 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  d2_5 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  d2_6 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  d2_7 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  d2_8 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  d2_9 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  d2_10 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  d2_11 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  d2_12 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  d2_13 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  d2_14 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  d2_15 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  d2_16 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  d2_17 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  d2_18 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  d2_19 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  d2_20 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  d2_21 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  d2_22 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  d2_23 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  d2_24 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  d2_25 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  d2_26 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  d2_27 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  d2_28 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  d2_29 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  d2_30 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  d2_31 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  age2_0 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  age2_1 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  age2_2 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  age2_3 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  age2_4 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  age2_5 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  age2_6 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  age2_7 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  age2_8 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  age2_9 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  age2_10 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  age2_11 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  age2_12 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  age2_13 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  age2_14 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  age2_15 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  age2_16 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  age2_17 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  age2_18 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  age2_19 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  age2_20 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  age2_21 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  age2_22 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  age2_23 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  age2_24 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  age2_25 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  age2_26 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  age2_27 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  age2_28 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  age2_29 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  age2_30 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  age2_31 = _RAND_259[0:0];
  _RAND_260 = {2{`RANDOM}};
  tag2_0 = _RAND_260[52:0];
  _RAND_261 = {2{`RANDOM}};
  tag2_1 = _RAND_261[52:0];
  _RAND_262 = {2{`RANDOM}};
  tag2_2 = _RAND_262[52:0];
  _RAND_263 = {2{`RANDOM}};
  tag2_3 = _RAND_263[52:0];
  _RAND_264 = {2{`RANDOM}};
  tag2_4 = _RAND_264[52:0];
  _RAND_265 = {2{`RANDOM}};
  tag2_5 = _RAND_265[52:0];
  _RAND_266 = {2{`RANDOM}};
  tag2_6 = _RAND_266[52:0];
  _RAND_267 = {2{`RANDOM}};
  tag2_7 = _RAND_267[52:0];
  _RAND_268 = {2{`RANDOM}};
  tag2_8 = _RAND_268[52:0];
  _RAND_269 = {2{`RANDOM}};
  tag2_9 = _RAND_269[52:0];
  _RAND_270 = {2{`RANDOM}};
  tag2_10 = _RAND_270[52:0];
  _RAND_271 = {2{`RANDOM}};
  tag2_11 = _RAND_271[52:0];
  _RAND_272 = {2{`RANDOM}};
  tag2_12 = _RAND_272[52:0];
  _RAND_273 = {2{`RANDOM}};
  tag2_13 = _RAND_273[52:0];
  _RAND_274 = {2{`RANDOM}};
  tag2_14 = _RAND_274[52:0];
  _RAND_275 = {2{`RANDOM}};
  tag2_15 = _RAND_275[52:0];
  _RAND_276 = {2{`RANDOM}};
  tag2_16 = _RAND_276[52:0];
  _RAND_277 = {2{`RANDOM}};
  tag2_17 = _RAND_277[52:0];
  _RAND_278 = {2{`RANDOM}};
  tag2_18 = _RAND_278[52:0];
  _RAND_279 = {2{`RANDOM}};
  tag2_19 = _RAND_279[52:0];
  _RAND_280 = {2{`RANDOM}};
  tag2_20 = _RAND_280[52:0];
  _RAND_281 = {2{`RANDOM}};
  tag2_21 = _RAND_281[52:0];
  _RAND_282 = {2{`RANDOM}};
  tag2_22 = _RAND_282[52:0];
  _RAND_283 = {2{`RANDOM}};
  tag2_23 = _RAND_283[52:0];
  _RAND_284 = {2{`RANDOM}};
  tag2_24 = _RAND_284[52:0];
  _RAND_285 = {2{`RANDOM}};
  tag2_25 = _RAND_285[52:0];
  _RAND_286 = {2{`RANDOM}};
  tag2_26 = _RAND_286[52:0];
  _RAND_287 = {2{`RANDOM}};
  tag2_27 = _RAND_287[52:0];
  _RAND_288 = {2{`RANDOM}};
  tag2_28 = _RAND_288[52:0];
  _RAND_289 = {2{`RANDOM}};
  tag2_29 = _RAND_289[52:0];
  _RAND_290 = {2{`RANDOM}};
  tag2_30 = _RAND_290[52:0];
  _RAND_291 = {2{`RANDOM}};
  tag2_31 = _RAND_291[52:0];
  _RAND_292 = {16{`RANDOM}};
  block2_0 = _RAND_292[511:0];
  _RAND_293 = {16{`RANDOM}};
  block2_1 = _RAND_293[511:0];
  _RAND_294 = {16{`RANDOM}};
  block2_2 = _RAND_294[511:0];
  _RAND_295 = {16{`RANDOM}};
  block2_3 = _RAND_295[511:0];
  _RAND_296 = {16{`RANDOM}};
  block2_4 = _RAND_296[511:0];
  _RAND_297 = {16{`RANDOM}};
  block2_5 = _RAND_297[511:0];
  _RAND_298 = {16{`RANDOM}};
  block2_6 = _RAND_298[511:0];
  _RAND_299 = {16{`RANDOM}};
  block2_7 = _RAND_299[511:0];
  _RAND_300 = {16{`RANDOM}};
  block2_8 = _RAND_300[511:0];
  _RAND_301 = {16{`RANDOM}};
  block2_9 = _RAND_301[511:0];
  _RAND_302 = {16{`RANDOM}};
  block2_10 = _RAND_302[511:0];
  _RAND_303 = {16{`RANDOM}};
  block2_11 = _RAND_303[511:0];
  _RAND_304 = {16{`RANDOM}};
  block2_12 = _RAND_304[511:0];
  _RAND_305 = {16{`RANDOM}};
  block2_13 = _RAND_305[511:0];
  _RAND_306 = {16{`RANDOM}};
  block2_14 = _RAND_306[511:0];
  _RAND_307 = {16{`RANDOM}};
  block2_15 = _RAND_307[511:0];
  _RAND_308 = {16{`RANDOM}};
  block2_16 = _RAND_308[511:0];
  _RAND_309 = {16{`RANDOM}};
  block2_17 = _RAND_309[511:0];
  _RAND_310 = {16{`RANDOM}};
  block2_18 = _RAND_310[511:0];
  _RAND_311 = {16{`RANDOM}};
  block2_19 = _RAND_311[511:0];
  _RAND_312 = {16{`RANDOM}};
  block2_20 = _RAND_312[511:0];
  _RAND_313 = {16{`RANDOM}};
  block2_21 = _RAND_313[511:0];
  _RAND_314 = {16{`RANDOM}};
  block2_22 = _RAND_314[511:0];
  _RAND_315 = {16{`RANDOM}};
  block2_23 = _RAND_315[511:0];
  _RAND_316 = {16{`RANDOM}};
  block2_24 = _RAND_316[511:0];
  _RAND_317 = {16{`RANDOM}};
  block2_25 = _RAND_317[511:0];
  _RAND_318 = {16{`RANDOM}};
  block2_26 = _RAND_318[511:0];
  _RAND_319 = {16{`RANDOM}};
  block2_27 = _RAND_319[511:0];
  _RAND_320 = {16{`RANDOM}};
  block2_28 = _RAND_320[511:0];
  _RAND_321 = {16{`RANDOM}};
  block2_29 = _RAND_321[511:0];
  _RAND_322 = {16{`RANDOM}};
  block2_30 = _RAND_322[511:0];
  _RAND_323 = {16{`RANDOM}};
  block2_31 = _RAND_323[511:0];
  _RAND_324 = {1{`RANDOM}};
  state = _RAND_324[1:0];
  _RAND_325 = {1{`RANDOM}};
  not_en_yet = _RAND_325[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI(
  input          clock,
  input          reset,
  input          io_out_aw_ready,
  output         io_out_aw_valid,
  output [63:0]  io_out_aw_bits_addr,
  input          io_out_w_ready,
  output         io_out_w_valid,
  output [63:0]  io_out_w_bits_data,
  output         io_out_w_bits_last,
  output         io_out_b_ready,
  input          io_out_b_valid,
  input          io_out_ar_ready,
  output         io_out_ar_valid,
  output [63:0]  io_out_ar_bits_addr,
  output         io_out_r_ready,
  input          io_out_r_valid,
  input  [63:0]  io_out_r_bits_data,
  input          io_out_r_bits_last,
  input          io_icacheio_req,
  input  [63:0]  io_icacheio_addr,
  output         io_icacheio_valid,
  output [511:0] io_icacheio_data,
  input          io_dcacheio_req,
  input  [63:0]  io_dcacheio_raddr,
  output         io_dcacheio_rvalid,
  output [511:0] io_dcacheio_rdata,
  input          io_dcacheio_weq,
  input  [63:0]  io_dcacheio_waddr,
  input  [511:0] io_dcacheio_wdata,
  output         io_dcacheio_wdone
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ibuffer_0; // @[AXI.scala 65:30]
  reg [63:0] ibuffer_1; // @[AXI.scala 65:30]
  reg [63:0] ibuffer_2; // @[AXI.scala 65:30]
  reg [63:0] ibuffer_3; // @[AXI.scala 65:30]
  reg [63:0] ibuffer_4; // @[AXI.scala 65:30]
  reg [63:0] ibuffer_5; // @[AXI.scala 65:30]
  reg [63:0] ibuffer_6; // @[AXI.scala 65:30]
  reg [63:0] ibuffer_7; // @[AXI.scala 65:30]
  reg [63:0] drbuffer_0; // @[AXI.scala 66:30]
  reg [63:0] drbuffer_1; // @[AXI.scala 66:30]
  reg [63:0] drbuffer_2; // @[AXI.scala 66:30]
  reg [63:0] drbuffer_3; // @[AXI.scala 66:30]
  reg [63:0] drbuffer_4; // @[AXI.scala 66:30]
  reg [63:0] drbuffer_5; // @[AXI.scala 66:30]
  reg [63:0] drbuffer_6; // @[AXI.scala 66:30]
  reg [63:0] drbuffer_7; // @[AXI.scala 66:30]
  reg [5:0] icnt; // @[AXI.scala 67:30]
  reg [5:0] drcnt; // @[AXI.scala 68:30]
  reg [5:0] dwcnt; // @[AXI.scala 69:30]
  reg [3:0] rstate; // @[AXI.scala 73:25]
  reg [2:0] wstate; // @[AXI.scala 74:25]
  wire  _T = 4'h0 == rstate; // @[Conditional.scala 37:30]
  wire  _T_1 = 4'h1 == rstate; // @[Conditional.scala 37:30]
  wire  _T_2 = 4'h2 == rstate; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_3 = io_out_r_valid ? 4'h3 : rstate; // @[AXI.scala 87:31 AXI.scala 87:39 AXI.scala 73:25]
  wire  _T_3 = 4'h3 == rstate; // @[Conditional.scala 37:30]
  wire  _T_5 = ~io_out_r_valid | io_out_r_bits_last; // @[AXI.scala 90:42]
  wire [3:0] _GEN_4 = ~io_out_r_valid | io_out_r_bits_last ? 4'h4 : rstate; // @[AXI.scala 90:62 AXI.scala 90:70 AXI.scala 73:25]
  wire  _T_6 = 4'h4 == rstate; // @[Conditional.scala 37:30]
  wire  _T_7 = 4'h5 == rstate; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_5 = io_out_ar_ready ? 4'h6 : rstate; // @[AXI.scala 97:32 AXI.scala 97:40 AXI.scala 73:25]
  wire  _T_8 = 4'h6 == rstate; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_6 = io_out_r_valid ? 4'h7 : rstate; // @[AXI.scala 100:31 AXI.scala 100:39 AXI.scala 73:25]
  wire  _T_9 = 4'h7 == rstate; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_7 = _T_5 ? 4'h8 : rstate; // @[AXI.scala 103:62 AXI.scala 103:70 AXI.scala 73:25]
  wire  _T_12 = 4'h8 == rstate; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_8 = _T_12 ? 4'h0 : rstate; // @[Conditional.scala 39:67 AXI.scala 106:20 AXI.scala 73:25]
  wire [3:0] _GEN_9 = _T_9 ? _GEN_7 : _GEN_8; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_10 = _T_8 ? _GEN_6 : _GEN_9; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_11 = _T_7 ? _GEN_5 : _GEN_10; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_12 = _T_6 ? 4'h0 : _GEN_11; // @[Conditional.scala 39:67 AXI.scala 93:20]
  wire [3:0] _GEN_13 = _T_3 ? _GEN_4 : _GEN_12; // @[Conditional.scala 39:67]
  wire  _T_13 = 3'h0 == wstate; // @[Conditional.scala 37:30]
  wire  _T_14 = 3'h1 == wstate; // @[Conditional.scala 37:30]
  wire  _T_15 = 3'h2 == wstate; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_19 = io_out_w_bits_last ? 3'h3 : wstate; // @[AXI.scala 119:35 AXI.scala 119:43 AXI.scala 74:25]
  wire  _T_16 = 3'h3 == wstate; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_20 = io_out_b_valid ? 3'h4 : wstate; // @[AXI.scala 122:31 AXI.scala 122:39 AXI.scala 74:25]
  wire  _T_17 = 3'h4 == wstate; // @[Conditional.scala 37:30]
  wire  _T_18 = ~io_out_b_valid; // @[AXI.scala 125:18]
  wire [2:0] _GEN_21 = ~io_out_b_valid ? 3'h0 : wstate; // @[AXI.scala 125:32 AXI.scala 125:40 AXI.scala 74:25]
  wire [2:0] _GEN_22 = _T_17 ? _GEN_21 : wstate; // @[Conditional.scala 39:67 AXI.scala 74:25]
  wire [2:0] _GEN_23 = _T_16 ? _GEN_20 : _GEN_22; // @[Conditional.scala 39:67]
  wire  _ibuffer_T = rstate == 4'h3; // @[AXI.scala 131:33]
  wire [63:0] _GEN_28 = 3'h1 == icnt[2:0] ? ibuffer_1 : ibuffer_0; // @[AXI.scala 131:25 AXI.scala 131:25]
  wire [63:0] _GEN_29 = 3'h2 == icnt[2:0] ? ibuffer_2 : _GEN_28; // @[AXI.scala 131:25 AXI.scala 131:25]
  wire [63:0] _GEN_30 = 3'h3 == icnt[2:0] ? ibuffer_3 : _GEN_29; // @[AXI.scala 131:25 AXI.scala 131:25]
  wire [63:0] _GEN_31 = 3'h4 == icnt[2:0] ? ibuffer_4 : _GEN_30; // @[AXI.scala 131:25 AXI.scala 131:25]
  wire [63:0] _GEN_32 = 3'h5 == icnt[2:0] ? ibuffer_5 : _GEN_31; // @[AXI.scala 131:25 AXI.scala 131:25]
  wire [63:0] _GEN_33 = 3'h6 == icnt[2:0] ? ibuffer_6 : _GEN_32; // @[AXI.scala 131:25 AXI.scala 131:25]
  wire [5:0] _icnt_T_2 = icnt + 6'h1; // @[AXI.scala 132:42]
  wire  _drbuffer_T = rstate == 4'h7; // @[AXI.scala 133:35]
  wire [63:0] _GEN_44 = 3'h1 == drcnt[2:0] ? drbuffer_1 : drbuffer_0; // @[AXI.scala 133:27 AXI.scala 133:27]
  wire [63:0] _GEN_45 = 3'h2 == drcnt[2:0] ? drbuffer_2 : _GEN_44; // @[AXI.scala 133:27 AXI.scala 133:27]
  wire [63:0] _GEN_46 = 3'h3 == drcnt[2:0] ? drbuffer_3 : _GEN_45; // @[AXI.scala 133:27 AXI.scala 133:27]
  wire [63:0] _GEN_47 = 3'h4 == drcnt[2:0] ? drbuffer_4 : _GEN_46; // @[AXI.scala 133:27 AXI.scala 133:27]
  wire [63:0] _GEN_48 = 3'h5 == drcnt[2:0] ? drbuffer_5 : _GEN_47; // @[AXI.scala 133:27 AXI.scala 133:27]
  wire [63:0] _GEN_49 = 3'h6 == drcnt[2:0] ? drbuffer_6 : _GEN_48; // @[AXI.scala 133:27 AXI.scala 133:27]
  wire [5:0] _drcnt_T_2 = drcnt + 6'h1; // @[AXI.scala 134:44]
  wire [5:0] _dwcnt_T_3 = dwcnt + 6'h1; // @[AXI.scala 135:58]
  wire [447:0] lo_5 = {ibuffer_6,ibuffer_5,ibuffer_4,ibuffer_3,ibuffer_2,ibuffer_1,ibuffer_0}; // @[Cat.scala 30:58]
  wire [447:0] lo_11 = {drbuffer_6,drbuffer_5,drbuffer_4,drbuffer_3,drbuffer_2,drbuffer_1,drbuffer_0}; // @[Cat.scala 30:58]
  wire  _io_out_ar_valid_T = rstate == 4'h1; // @[AXI.scala 160:35]
  wire  _io_out_ar_valid_T_1 = rstate == 4'h5; // @[AXI.scala 160:57]
  wire [63:0] _io_out_ar_bits_addr_T_2 = _io_out_ar_valid_T_1 ? io_dcacheio_raddr : 64'h0; // @[AXI.scala 161:70]
  wire [11:0] _io_out_w_bits_data_T = {dwcnt, 6'h0}; // @[AXI.scala 196:54]
  wire [511:0] _io_out_w_bits_data_T_1 = io_dcacheio_wdata >> _io_out_w_bits_data_T; // @[AXI.scala 196:44]
  assign io_out_aw_valid = wstate == 3'h1; // @[AXI.scala 183:35]
  assign io_out_aw_bits_addr = io_dcacheio_waddr; // @[AXI.scala 184:25]
  assign io_out_w_valid = wstate == 3'h2; // @[AXI.scala 195:35]
  assign io_out_w_bits_data = _io_out_w_bits_data_T_1[63:0]; // @[AXI.scala 196:60]
  assign io_out_w_bits_last = dwcnt == 6'h8; // @[AXI.scala 198:34]
  assign io_out_b_ready = wstate == 3'h4; // @[AXI.scala 200:35]
  assign io_out_ar_valid = rstate == 4'h1 | rstate == 4'h5; // @[AXI.scala 160:47]
  assign io_out_ar_bits_addr = _io_out_ar_valid_T ? io_icacheio_addr : _io_out_ar_bits_addr_T_2; // @[AXI.scala 161:31]
  assign io_out_r_ready = _ibuffer_T | _drbuffer_T; // @[AXI.scala 179:47]
  assign io_icacheio_valid = rstate == 4'h4; // @[AXI.scala 144:31]
  assign io_icacheio_data = {ibuffer_7,lo_5}; // @[Cat.scala 30:58]
  assign io_dcacheio_rvalid = rstate == 4'h8; // @[AXI.scala 151:31]
  assign io_dcacheio_rdata = {drbuffer_7,lo_11}; // @[Cat.scala 30:58]
  assign io_dcacheio_wdone = wstate == 3'h4 & _T_18; // @[AXI.scala 154:42]
  always @(posedge clock) begin
    if (reset) begin // @[AXI.scala 65:30]
      ibuffer_0 <= 64'h0; // @[AXI.scala 65:30]
    end else if (3'h0 == icnt[2:0]) begin // @[AXI.scala 131:19]
      if (rstate == 4'h3) begin // @[AXI.scala 131:25]
        ibuffer_0 <= io_out_r_bits_data;
      end else if (3'h7 == icnt[2:0]) begin // @[AXI.scala 131:25]
        ibuffer_0 <= ibuffer_7; // @[AXI.scala 131:25]
      end else begin
        ibuffer_0 <= _GEN_33;
      end
    end
    if (reset) begin // @[AXI.scala 65:30]
      ibuffer_1 <= 64'h0; // @[AXI.scala 65:30]
    end else if (3'h1 == icnt[2:0]) begin // @[AXI.scala 131:19]
      if (rstate == 4'h3) begin // @[AXI.scala 131:25]
        ibuffer_1 <= io_out_r_bits_data;
      end else if (3'h7 == icnt[2:0]) begin // @[AXI.scala 131:25]
        ibuffer_1 <= ibuffer_7; // @[AXI.scala 131:25]
      end else begin
        ibuffer_1 <= _GEN_33;
      end
    end
    if (reset) begin // @[AXI.scala 65:30]
      ibuffer_2 <= 64'h0; // @[AXI.scala 65:30]
    end else if (3'h2 == icnt[2:0]) begin // @[AXI.scala 131:19]
      if (rstate == 4'h3) begin // @[AXI.scala 131:25]
        ibuffer_2 <= io_out_r_bits_data;
      end else if (3'h7 == icnt[2:0]) begin // @[AXI.scala 131:25]
        ibuffer_2 <= ibuffer_7; // @[AXI.scala 131:25]
      end else begin
        ibuffer_2 <= _GEN_33;
      end
    end
    if (reset) begin // @[AXI.scala 65:30]
      ibuffer_3 <= 64'h0; // @[AXI.scala 65:30]
    end else if (3'h3 == icnt[2:0]) begin // @[AXI.scala 131:19]
      if (rstate == 4'h3) begin // @[AXI.scala 131:25]
        ibuffer_3 <= io_out_r_bits_data;
      end else if (3'h7 == icnt[2:0]) begin // @[AXI.scala 131:25]
        ibuffer_3 <= ibuffer_7; // @[AXI.scala 131:25]
      end else begin
        ibuffer_3 <= _GEN_33;
      end
    end
    if (reset) begin // @[AXI.scala 65:30]
      ibuffer_4 <= 64'h0; // @[AXI.scala 65:30]
    end else if (3'h4 == icnt[2:0]) begin // @[AXI.scala 131:19]
      if (rstate == 4'h3) begin // @[AXI.scala 131:25]
        ibuffer_4 <= io_out_r_bits_data;
      end else if (3'h7 == icnt[2:0]) begin // @[AXI.scala 131:25]
        ibuffer_4 <= ibuffer_7; // @[AXI.scala 131:25]
      end else begin
        ibuffer_4 <= _GEN_33;
      end
    end
    if (reset) begin // @[AXI.scala 65:30]
      ibuffer_5 <= 64'h0; // @[AXI.scala 65:30]
    end else if (3'h5 == icnt[2:0]) begin // @[AXI.scala 131:19]
      if (rstate == 4'h3) begin // @[AXI.scala 131:25]
        ibuffer_5 <= io_out_r_bits_data;
      end else if (3'h7 == icnt[2:0]) begin // @[AXI.scala 131:25]
        ibuffer_5 <= ibuffer_7; // @[AXI.scala 131:25]
      end else begin
        ibuffer_5 <= _GEN_33;
      end
    end
    if (reset) begin // @[AXI.scala 65:30]
      ibuffer_6 <= 64'h0; // @[AXI.scala 65:30]
    end else if (3'h6 == icnt[2:0]) begin // @[AXI.scala 131:19]
      if (rstate == 4'h3) begin // @[AXI.scala 131:25]
        ibuffer_6 <= io_out_r_bits_data;
      end else if (3'h7 == icnt[2:0]) begin // @[AXI.scala 131:25]
        ibuffer_6 <= ibuffer_7; // @[AXI.scala 131:25]
      end else begin
        ibuffer_6 <= _GEN_33;
      end
    end
    if (reset) begin // @[AXI.scala 65:30]
      ibuffer_7 <= 64'h0; // @[AXI.scala 65:30]
    end else if (3'h7 == icnt[2:0]) begin // @[AXI.scala 131:19]
      if (rstate == 4'h3) begin // @[AXI.scala 131:25]
        ibuffer_7 <= io_out_r_bits_data;
      end else if (!(3'h7 == icnt[2:0])) begin // @[AXI.scala 131:25]
        ibuffer_7 <= _GEN_33;
      end
    end
    if (reset) begin // @[AXI.scala 66:30]
      drbuffer_0 <= 64'h0; // @[AXI.scala 66:30]
    end else if (3'h0 == drcnt[2:0]) begin // @[AXI.scala 133:21]
      if (rstate == 4'h7) begin // @[AXI.scala 133:27]
        drbuffer_0 <= io_out_r_bits_data;
      end else if (3'h7 == drcnt[2:0]) begin // @[AXI.scala 133:27]
        drbuffer_0 <= drbuffer_7; // @[AXI.scala 133:27]
      end else begin
        drbuffer_0 <= _GEN_49;
      end
    end
    if (reset) begin // @[AXI.scala 66:30]
      drbuffer_1 <= 64'h0; // @[AXI.scala 66:30]
    end else if (3'h1 == drcnt[2:0]) begin // @[AXI.scala 133:21]
      if (rstate == 4'h7) begin // @[AXI.scala 133:27]
        drbuffer_1 <= io_out_r_bits_data;
      end else if (3'h7 == drcnt[2:0]) begin // @[AXI.scala 133:27]
        drbuffer_1 <= drbuffer_7; // @[AXI.scala 133:27]
      end else begin
        drbuffer_1 <= _GEN_49;
      end
    end
    if (reset) begin // @[AXI.scala 66:30]
      drbuffer_2 <= 64'h0; // @[AXI.scala 66:30]
    end else if (3'h2 == drcnt[2:0]) begin // @[AXI.scala 133:21]
      if (rstate == 4'h7) begin // @[AXI.scala 133:27]
        drbuffer_2 <= io_out_r_bits_data;
      end else if (3'h7 == drcnt[2:0]) begin // @[AXI.scala 133:27]
        drbuffer_2 <= drbuffer_7; // @[AXI.scala 133:27]
      end else begin
        drbuffer_2 <= _GEN_49;
      end
    end
    if (reset) begin // @[AXI.scala 66:30]
      drbuffer_3 <= 64'h0; // @[AXI.scala 66:30]
    end else if (3'h3 == drcnt[2:0]) begin // @[AXI.scala 133:21]
      if (rstate == 4'h7) begin // @[AXI.scala 133:27]
        drbuffer_3 <= io_out_r_bits_data;
      end else if (3'h7 == drcnt[2:0]) begin // @[AXI.scala 133:27]
        drbuffer_3 <= drbuffer_7; // @[AXI.scala 133:27]
      end else begin
        drbuffer_3 <= _GEN_49;
      end
    end
    if (reset) begin // @[AXI.scala 66:30]
      drbuffer_4 <= 64'h0; // @[AXI.scala 66:30]
    end else if (3'h4 == drcnt[2:0]) begin // @[AXI.scala 133:21]
      if (rstate == 4'h7) begin // @[AXI.scala 133:27]
        drbuffer_4 <= io_out_r_bits_data;
      end else if (3'h7 == drcnt[2:0]) begin // @[AXI.scala 133:27]
        drbuffer_4 <= drbuffer_7; // @[AXI.scala 133:27]
      end else begin
        drbuffer_4 <= _GEN_49;
      end
    end
    if (reset) begin // @[AXI.scala 66:30]
      drbuffer_5 <= 64'h0; // @[AXI.scala 66:30]
    end else if (3'h5 == drcnt[2:0]) begin // @[AXI.scala 133:21]
      if (rstate == 4'h7) begin // @[AXI.scala 133:27]
        drbuffer_5 <= io_out_r_bits_data;
      end else if (3'h7 == drcnt[2:0]) begin // @[AXI.scala 133:27]
        drbuffer_5 <= drbuffer_7; // @[AXI.scala 133:27]
      end else begin
        drbuffer_5 <= _GEN_49;
      end
    end
    if (reset) begin // @[AXI.scala 66:30]
      drbuffer_6 <= 64'h0; // @[AXI.scala 66:30]
    end else if (3'h6 == drcnt[2:0]) begin // @[AXI.scala 133:21]
      if (rstate == 4'h7) begin // @[AXI.scala 133:27]
        drbuffer_6 <= io_out_r_bits_data;
      end else if (3'h7 == drcnt[2:0]) begin // @[AXI.scala 133:27]
        drbuffer_6 <= drbuffer_7; // @[AXI.scala 133:27]
      end else begin
        drbuffer_6 <= _GEN_49;
      end
    end
    if (reset) begin // @[AXI.scala 66:30]
      drbuffer_7 <= 64'h0; // @[AXI.scala 66:30]
    end else if (3'h7 == drcnt[2:0]) begin // @[AXI.scala 133:21]
      if (rstate == 4'h7) begin // @[AXI.scala 133:27]
        drbuffer_7 <= io_out_r_bits_data;
      end else if (!(3'h7 == drcnt[2:0])) begin // @[AXI.scala 133:27]
        drbuffer_7 <= _GEN_49;
      end
    end
    if (reset) begin // @[AXI.scala 67:30]
      icnt <= 6'h0; // @[AXI.scala 67:30]
    end else if (_ibuffer_T) begin // @[AXI.scala 132:16]
      icnt <= _icnt_T_2;
    end else begin
      icnt <= 6'h0;
    end
    if (reset) begin // @[AXI.scala 68:30]
      drcnt <= 6'h0; // @[AXI.scala 68:30]
    end else if (_drbuffer_T) begin // @[AXI.scala 134:17]
      drcnt <= _drcnt_T_2;
    end else begin
      drcnt <= 6'h0;
    end
    if (reset) begin // @[AXI.scala 69:30]
      dwcnt <= 6'h0; // @[AXI.scala 69:30]
    end else if (wstate == 3'h2 & io_out_w_ready) begin // @[AXI.scala 135:17]
      dwcnt <= _dwcnt_T_3;
    end else begin
      dwcnt <= 6'h0;
    end
    if (reset) begin // @[AXI.scala 73:25]
      rstate <= 4'h0; // @[AXI.scala 73:25]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_icacheio_req) begin // @[AXI.scala 79:32]
        rstate <= 4'h1; // @[AXI.scala 79:40]
      end else if (io_dcacheio_req) begin // @[AXI.scala 80:37]
        rstate <= 4'h5; // @[AXI.scala 80:45]
      end
    end else if (_T_1) begin // @[Conditional.scala 39:67]
      if (io_out_ar_ready) begin // @[AXI.scala 84:32]
        rstate <= 4'h2; // @[AXI.scala 84:40]
      end
    end else if (_T_2) begin // @[Conditional.scala 39:67]
      rstate <= _GEN_3;
    end else begin
      rstate <= _GEN_13;
    end
    if (reset) begin // @[AXI.scala 74:25]
      wstate <= 3'h0; // @[AXI.scala 74:25]
    end else if (_T_13) begin // @[Conditional.scala 40:58]
      if (io_dcacheio_weq) begin // @[AXI.scala 113:32]
        wstate <= 3'h1; // @[AXI.scala 113:40]
      end
    end else if (_T_14) begin // @[Conditional.scala 39:67]
      if (io_out_aw_ready) begin // @[AXI.scala 116:32]
        wstate <= 3'h2; // @[AXI.scala 116:40]
      end
    end else if (_T_15) begin // @[Conditional.scala 39:67]
      wstate <= _GEN_19;
    end else begin
      wstate <= _GEN_23;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  ibuffer_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  ibuffer_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  ibuffer_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  ibuffer_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  ibuffer_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  ibuffer_5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  ibuffer_6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  ibuffer_7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  drbuffer_0 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  drbuffer_1 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  drbuffer_2 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  drbuffer_3 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  drbuffer_4 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  drbuffer_5 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  drbuffer_6 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  drbuffer_7 = _RAND_15[63:0];
  _RAND_16 = {1{`RANDOM}};
  icnt = _RAND_16[5:0];
  _RAND_17 = {1{`RANDOM}};
  drcnt = _RAND_17[5:0];
  _RAND_18 = {1{`RANDOM}};
  dwcnt = _RAND_18[5:0];
  _RAND_19 = {1{`RANDOM}};
  rstate = _RAND_19[3:0];
  _RAND_20 = {1{`RANDOM}};
  wstate = _RAND_20[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Clint(
  input         clock,
  input         reset,
  input         io_dmem_en,
  input         io_dmem_op,
  input  [63:0] io_dmem_addr,
  input  [63:0] io_dmem_wdata,
  input  [7:0]  io_dmem_wmask,
  output        io_dmem_ok,
  output [63:0] io_dmem_rdata,
  output        io_mem0_en,
  output        io_mem0_op,
  output [63:0] io_mem0_addr,
  output [63:0] io_mem0_wdata,
  output [7:0]  io_mem0_wmask,
  input         io_mem0_ok,
  input  [63:0] io_mem0_rdata,
  input  [63:0] io_mem1_rdata,
  output        io_mem2_en,
  output        io_mem2_op,
  output [63:0] io_mem2_wdata,
  output [7:0]  io_mem2_wmask,
  input  [63:0] io_mem2_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [1:0] _GEN_0 = io_dmem_addr == 64'h2004000 ? 2'h2 : 2'h0; // @[Clint.scala 21:50 Clint.scala 21:55 Clint.scala 22:24]
  wire [1:0] _GEN_1 = io_dmem_addr == 64'h200bff8 ? 2'h1 : _GEN_0; // @[Clint.scala 20:45 Clint.scala 20:50]
  wire [1:0] sel = ~io_mem0_ok ? 2'h0 : _GEN_1; // @[Clint.scala 16:22 Clint.scala 16:27]
  reg [1:0] sel_r; // @[Reg.scala 27:20]
  wire  out_ok = 2'h2 == sel_r | (2'h1 == sel_r | 2'h0 == sel_r & io_mem0_ok); // @[Mux.scala 80:57]
  wire  _io_mem0_en_T = sel == 2'h0; // @[Clint.scala 27:32]
  wire  _io_mem2_en_T = sel == 2'h2; // @[Clint.scala 37:32]
  wire [63:0] _out_rdata_T_1 = 2'h0 == sel_r ? io_mem0_rdata : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _out_rdata_T_3 = 2'h1 == sel_r ? io_mem1_rdata : _out_rdata_T_1; // @[Mux.scala 80:57]
  assign io_dmem_ok = 2'h2 == sel_r | (2'h1 == sel_r | 2'h0 == sel_r & io_mem0_ok); // @[Mux.scala 80:57]
  assign io_dmem_rdata = 2'h2 == sel_r ? io_mem2_rdata : _out_rdata_T_3; // @[Mux.scala 80:57]
  assign io_mem0_en = sel == 2'h0 & io_dmem_en; // @[Clint.scala 27:27]
  assign io_mem0_op = _io_mem0_en_T & io_dmem_op; // @[Clint.scala 28:27]
  assign io_mem0_addr = _io_mem0_en_T ? io_dmem_addr : 64'h0; // @[Clint.scala 29:27]
  assign io_mem0_wdata = _io_mem0_en_T ? io_dmem_wdata : 64'h0; // @[Clint.scala 30:27]
  assign io_mem0_wmask = _io_mem0_en_T ? io_dmem_wmask : 8'h0; // @[Clint.scala 31:27]
  assign io_mem2_en = sel == 2'h2 & io_dmem_en; // @[Clint.scala 37:27]
  assign io_mem2_op = _io_mem2_en_T & io_dmem_op; // @[Clint.scala 38:27]
  assign io_mem2_wdata = _io_mem2_en_T ? io_dmem_wdata : 64'h0; // @[Clint.scala 40:27]
  assign io_mem2_wmask = _io_mem2_en_T ? io_dmem_wmask : 8'h0; // @[Clint.scala 41:27]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 27:20]
      sel_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (out_ok) begin // @[Reg.scala 28:19]
      if (~io_mem0_ok) begin // @[Clint.scala 16:22]
        sel_r <= 2'h0; // @[Clint.scala 16:27]
      end else if (io_dmem_addr == 64'h200bff8) begin // @[Clint.scala 20:45]
        sel_r <= 2'h1; // @[Clint.scala 20:50]
      end else begin
        sel_r <= _GEN_0;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sel_r = _RAND_0[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Mtime(
  input         clock,
  input         reset,
  output [63:0] io_mem_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] mtime; // @[Clint.scala 63:24]
  wire [63:0] _mtime_T_1 = mtime + 64'h1; // @[Clint.scala 64:20]
  assign io_mem_rdata = mtime; // @[Clint.scala 67:18]
  always @(posedge clock) begin
    if (reset) begin // @[Clint.scala 63:24]
      mtime <= 64'h0; // @[Clint.scala 63:24]
    end else begin
      mtime <= _mtime_T_1; // @[Clint.scala 64:11]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mtime = _RAND_0[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Mtimecmp(
  input         clock,
  input         reset,
  input         io_mem_en,
  input         io_mem_op,
  input  [63:0] io_mem_wdata,
  input  [7:0]  io_mem_wmask,
  output [63:0] io_mem_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] mtimecmp; // @[Clint.scala 74:27]
  wire [7:0] mask64_hi_hi_hi = io_mem_wmask[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] mask64_hi_hi_lo = io_mem_wmask[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] mask64_hi_lo_hi = io_mem_wmask[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] mask64_hi_lo_lo = io_mem_wmask[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] mask64_lo_hi_hi = io_mem_wmask[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] mask64_lo_hi_lo = io_mem_wmask[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] mask64_lo_lo_hi = io_mem_wmask[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] mask64_lo_lo_lo = io_mem_wmask[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [63:0] mask64 = {mask64_hi_hi_hi,mask64_hi_hi_lo,mask64_hi_lo_hi,mask64_hi_lo_lo,mask64_lo_hi_hi,mask64_lo_hi_lo,
    mask64_lo_lo_hi,mask64_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [63:0] _mtimecmp_update_T = ~mask64; // @[Clint.scala 78:40]
  wire [63:0] _mtimecmp_update_T_1 = mtimecmp & _mtimecmp_update_T; // @[Clint.scala 78:37]
  wire [63:0] _mtimecmp_update_T_2 = mask64 & io_mem_wdata; // @[Clint.scala 78:60]
  wire [63:0] mtimecmp_update = _mtimecmp_update_T_1 | _mtimecmp_update_T_2; // @[Clint.scala 78:50]
  assign io_mem_rdata = mtimecmp; // @[Clint.scala 83:18]
  always @(posedge clock) begin
    if (reset) begin // @[Clint.scala 74:27]
      mtimecmp <= 64'h0; // @[Clint.scala 74:27]
    end else if (io_mem_en & io_mem_op) begin // @[Clint.scala 80:33]
      mtimecmp <= mtimecmp_update; // @[Clint.scala 80:43]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mtimecmp = _RAND_0[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SimTop(
  input         clock,
  input         reset,
  input  [63:0] io_logCtrl_log_begin,
  input  [63:0] io_logCtrl_log_end,
  input  [63:0] io_logCtrl_log_level,
  input         io_perfInfo_clean,
  input         io_perfInfo_dump,
  output        io_uart_out_valid,
  output [7:0]  io_uart_out_ch,
  output        io_uart_in_valid,
  input  [7:0]  io_uart_in_ch,
  input         io_memAXI_0_aw_ready,
  output        io_memAXI_0_aw_valid,
  output [7:0]  io_memAXI_0_aw_bits_len,
  output [2:0]  io_memAXI_0_aw_bits_size,
  output [1:0]  io_memAXI_0_aw_bits_burst,
  output        io_memAXI_0_aw_bits_lock,
  output [3:0]  io_memAXI_0_aw_bits_cache,
  output [3:0]  io_memAXI_0_aw_bits_qos,
  output [63:0] io_memAXI_0_aw_bits_addr,
  output [2:0]  io_memAXI_0_aw_bits_prot,
  output [3:0]  io_memAXI_0_aw_bits_id,
  output [3:0]  io_memAXI_0_aw_bits_user,
  input         io_memAXI_0_w_ready,
  output        io_memAXI_0_w_valid,
  output [63:0] io_memAXI_0_w_bits_data,
  output [7:0]  io_memAXI_0_w_bits_strb,
  output        io_memAXI_0_w_bits_last,
  output        io_memAXI_0_b_ready,
  input         io_memAXI_0_b_valid,
  input  [1:0]  io_memAXI_0_b_bits_resp,
  input  [3:0]  io_memAXI_0_b_bits_id,
  input  [3:0]  io_memAXI_0_b_bits_user,
  input         io_memAXI_0_ar_ready,
  output        io_memAXI_0_ar_valid,
  output [7:0]  io_memAXI_0_ar_bits_len,
  output [2:0]  io_memAXI_0_ar_bits_size,
  output [1:0]  io_memAXI_0_ar_bits_burst,
  output        io_memAXI_0_ar_bits_lock,
  output [3:0]  io_memAXI_0_ar_bits_cache,
  output [3:0]  io_memAXI_0_ar_bits_qos,
  output [63:0] io_memAXI_0_ar_bits_addr,
  output [2:0]  io_memAXI_0_ar_bits_prot,
  output [3:0]  io_memAXI_0_ar_bits_id,
  output [3:0]  io_memAXI_0_ar_bits_user,
  output        io_memAXI_0_r_ready,
  input         io_memAXI_0_r_valid,
  input  [1:0]  io_memAXI_0_r_bits_resp,
  input  [63:0] io_memAXI_0_r_bits_data,
  input         io_memAXI_0_r_bits_last,
  input  [3:0]  io_memAXI_0_r_bits_id,
  input  [3:0]  io_memAXI_0_r_bits_user
);
  wire  core_clock; // @[SimTop.scala 15:20]
  wire  core_reset; // @[SimTop.scala 15:20]
  wire [63:0] core_io_imem_addr; // @[SimTop.scala 15:20]
  wire [31:0] core_io_imem_data; // @[SimTop.scala 15:20]
  wire  core_io_imem_data_ok; // @[SimTop.scala 15:20]
  wire  core_io_dmem_en; // @[SimTop.scala 15:20]
  wire  core_io_dmem_op; // @[SimTop.scala 15:20]
  wire [63:0] core_io_dmem_addr; // @[SimTop.scala 15:20]
  wire [63:0] core_io_dmem_wdata; // @[SimTop.scala 15:20]
  wire [7:0] core_io_dmem_wmask; // @[SimTop.scala 15:20]
  wire  core_io_dmem_ok; // @[SimTop.scala 15:20]
  wire [63:0] core_io_dmem_rdata; // @[SimTop.scala 15:20]
  wire  icache_clock; // @[SimTop.scala 16:22]
  wire  icache_reset; // @[SimTop.scala 16:22]
  wire [63:0] icache_io_imem_addr; // @[SimTop.scala 16:22]
  wire [31:0] icache_io_imem_data; // @[SimTop.scala 16:22]
  wire  icache_io_imem_data_ok; // @[SimTop.scala 16:22]
  wire  icache_io_axi_req; // @[SimTop.scala 16:22]
  wire [63:0] icache_io_axi_addr; // @[SimTop.scala 16:22]
  wire  icache_io_axi_valid; // @[SimTop.scala 16:22]
  wire [511:0] icache_io_axi_data; // @[SimTop.scala 16:22]
  wire  dcache_clock; // @[SimTop.scala 17:22]
  wire  dcache_reset; // @[SimTop.scala 17:22]
  wire  dcache_io_dmem_en; // @[SimTop.scala 17:22]
  wire  dcache_io_dmem_op; // @[SimTop.scala 17:22]
  wire [63:0] dcache_io_dmem_addr; // @[SimTop.scala 17:22]
  wire [63:0] dcache_io_dmem_wdata; // @[SimTop.scala 17:22]
  wire [7:0] dcache_io_dmem_wmask; // @[SimTop.scala 17:22]
  wire  dcache_io_dmem_ok; // @[SimTop.scala 17:22]
  wire [63:0] dcache_io_dmem_rdata; // @[SimTop.scala 17:22]
  wire  dcache_io_axi_req; // @[SimTop.scala 17:22]
  wire [63:0] dcache_io_axi_raddr; // @[SimTop.scala 17:22]
  wire  dcache_io_axi_rvalid; // @[SimTop.scala 17:22]
  wire [511:0] dcache_io_axi_rdata; // @[SimTop.scala 17:22]
  wire  dcache_io_axi_weq; // @[SimTop.scala 17:22]
  wire [63:0] dcache_io_axi_waddr; // @[SimTop.scala 17:22]
  wire [511:0] dcache_io_axi_wdata; // @[SimTop.scala 17:22]
  wire  dcache_io_axi_wdone; // @[SimTop.scala 17:22]
  wire  axi_clock; // @[SimTop.scala 18:19]
  wire  axi_reset; // @[SimTop.scala 18:19]
  wire  axi_io_out_aw_ready; // @[SimTop.scala 18:19]
  wire  axi_io_out_aw_valid; // @[SimTop.scala 18:19]
  wire [63:0] axi_io_out_aw_bits_addr; // @[SimTop.scala 18:19]
  wire  axi_io_out_w_ready; // @[SimTop.scala 18:19]
  wire  axi_io_out_w_valid; // @[SimTop.scala 18:19]
  wire [63:0] axi_io_out_w_bits_data; // @[SimTop.scala 18:19]
  wire  axi_io_out_w_bits_last; // @[SimTop.scala 18:19]
  wire  axi_io_out_b_ready; // @[SimTop.scala 18:19]
  wire  axi_io_out_b_valid; // @[SimTop.scala 18:19]
  wire  axi_io_out_ar_ready; // @[SimTop.scala 18:19]
  wire  axi_io_out_ar_valid; // @[SimTop.scala 18:19]
  wire [63:0] axi_io_out_ar_bits_addr; // @[SimTop.scala 18:19]
  wire  axi_io_out_r_ready; // @[SimTop.scala 18:19]
  wire  axi_io_out_r_valid; // @[SimTop.scala 18:19]
  wire [63:0] axi_io_out_r_bits_data; // @[SimTop.scala 18:19]
  wire  axi_io_out_r_bits_last; // @[SimTop.scala 18:19]
  wire  axi_io_icacheio_req; // @[SimTop.scala 18:19]
  wire [63:0] axi_io_icacheio_addr; // @[SimTop.scala 18:19]
  wire  axi_io_icacheio_valid; // @[SimTop.scala 18:19]
  wire [511:0] axi_io_icacheio_data; // @[SimTop.scala 18:19]
  wire  axi_io_dcacheio_req; // @[SimTop.scala 18:19]
  wire [63:0] axi_io_dcacheio_raddr; // @[SimTop.scala 18:19]
  wire  axi_io_dcacheio_rvalid; // @[SimTop.scala 18:19]
  wire [511:0] axi_io_dcacheio_rdata; // @[SimTop.scala 18:19]
  wire  axi_io_dcacheio_weq; // @[SimTop.scala 18:19]
  wire [63:0] axi_io_dcacheio_waddr; // @[SimTop.scala 18:19]
  wire [511:0] axi_io_dcacheio_wdata; // @[SimTop.scala 18:19]
  wire  axi_io_dcacheio_wdone; // @[SimTop.scala 18:19]
  wire  clint_clock; // @[SimTop.scala 20:21]
  wire  clint_reset; // @[SimTop.scala 20:21]
  wire  clint_io_dmem_en; // @[SimTop.scala 20:21]
  wire  clint_io_dmem_op; // @[SimTop.scala 20:21]
  wire [63:0] clint_io_dmem_addr; // @[SimTop.scala 20:21]
  wire [63:0] clint_io_dmem_wdata; // @[SimTop.scala 20:21]
  wire [7:0] clint_io_dmem_wmask; // @[SimTop.scala 20:21]
  wire  clint_io_dmem_ok; // @[SimTop.scala 20:21]
  wire [63:0] clint_io_dmem_rdata; // @[SimTop.scala 20:21]
  wire  clint_io_mem0_en; // @[SimTop.scala 20:21]
  wire  clint_io_mem0_op; // @[SimTop.scala 20:21]
  wire [63:0] clint_io_mem0_addr; // @[SimTop.scala 20:21]
  wire [63:0] clint_io_mem0_wdata; // @[SimTop.scala 20:21]
  wire [7:0] clint_io_mem0_wmask; // @[SimTop.scala 20:21]
  wire  clint_io_mem0_ok; // @[SimTop.scala 20:21]
  wire [63:0] clint_io_mem0_rdata; // @[SimTop.scala 20:21]
  wire [63:0] clint_io_mem1_rdata; // @[SimTop.scala 20:21]
  wire  clint_io_mem2_en; // @[SimTop.scala 20:21]
  wire  clint_io_mem2_op; // @[SimTop.scala 20:21]
  wire [63:0] clint_io_mem2_wdata; // @[SimTop.scala 20:21]
  wire [7:0] clint_io_mem2_wmask; // @[SimTop.scala 20:21]
  wire [63:0] clint_io_mem2_rdata; // @[SimTop.scala 20:21]
  wire  mtime_clock; // @[SimTop.scala 21:21]
  wire  mtime_reset; // @[SimTop.scala 21:21]
  wire [63:0] mtime_io_mem_rdata; // @[SimTop.scala 21:21]
  wire  mtimecmp_clock; // @[SimTop.scala 22:24]
  wire  mtimecmp_reset; // @[SimTop.scala 22:24]
  wire  mtimecmp_io_mem_en; // @[SimTop.scala 22:24]
  wire  mtimecmp_io_mem_op; // @[SimTop.scala 22:24]
  wire [63:0] mtimecmp_io_mem_wdata; // @[SimTop.scala 22:24]
  wire [7:0] mtimecmp_io_mem_wmask; // @[SimTop.scala 22:24]
  wire [63:0] mtimecmp_io_mem_rdata; // @[SimTop.scala 22:24]
  Core core ( // @[SimTop.scala 15:20]
    .clock(core_clock),
    .reset(core_reset),
    .io_imem_addr(core_io_imem_addr),
    .io_imem_data(core_io_imem_data),
    .io_imem_data_ok(core_io_imem_data_ok),
    .io_dmem_en(core_io_dmem_en),
    .io_dmem_op(core_io_dmem_op),
    .io_dmem_addr(core_io_dmem_addr),
    .io_dmem_wdata(core_io_dmem_wdata),
    .io_dmem_wmask(core_io_dmem_wmask),
    .io_dmem_ok(core_io_dmem_ok),
    .io_dmem_rdata(core_io_dmem_rdata)
  );
  ICache icache ( // @[SimTop.scala 16:22]
    .clock(icache_clock),
    .reset(icache_reset),
    .io_imem_addr(icache_io_imem_addr),
    .io_imem_data(icache_io_imem_data),
    .io_imem_data_ok(icache_io_imem_data_ok),
    .io_axi_req(icache_io_axi_req),
    .io_axi_addr(icache_io_axi_addr),
    .io_axi_valid(icache_io_axi_valid),
    .io_axi_data(icache_io_axi_data)
  );
  DCache dcache ( // @[SimTop.scala 17:22]
    .clock(dcache_clock),
    .reset(dcache_reset),
    .io_dmem_en(dcache_io_dmem_en),
    .io_dmem_op(dcache_io_dmem_op),
    .io_dmem_addr(dcache_io_dmem_addr),
    .io_dmem_wdata(dcache_io_dmem_wdata),
    .io_dmem_wmask(dcache_io_dmem_wmask),
    .io_dmem_ok(dcache_io_dmem_ok),
    .io_dmem_rdata(dcache_io_dmem_rdata),
    .io_axi_req(dcache_io_axi_req),
    .io_axi_raddr(dcache_io_axi_raddr),
    .io_axi_rvalid(dcache_io_axi_rvalid),
    .io_axi_rdata(dcache_io_axi_rdata),
    .io_axi_weq(dcache_io_axi_weq),
    .io_axi_waddr(dcache_io_axi_waddr),
    .io_axi_wdata(dcache_io_axi_wdata),
    .io_axi_wdone(dcache_io_axi_wdone)
  );
  AXI axi ( // @[SimTop.scala 18:19]
    .clock(axi_clock),
    .reset(axi_reset),
    .io_out_aw_ready(axi_io_out_aw_ready),
    .io_out_aw_valid(axi_io_out_aw_valid),
    .io_out_aw_bits_addr(axi_io_out_aw_bits_addr),
    .io_out_w_ready(axi_io_out_w_ready),
    .io_out_w_valid(axi_io_out_w_valid),
    .io_out_w_bits_data(axi_io_out_w_bits_data),
    .io_out_w_bits_last(axi_io_out_w_bits_last),
    .io_out_b_ready(axi_io_out_b_ready),
    .io_out_b_valid(axi_io_out_b_valid),
    .io_out_ar_ready(axi_io_out_ar_ready),
    .io_out_ar_valid(axi_io_out_ar_valid),
    .io_out_ar_bits_addr(axi_io_out_ar_bits_addr),
    .io_out_r_ready(axi_io_out_r_ready),
    .io_out_r_valid(axi_io_out_r_valid),
    .io_out_r_bits_data(axi_io_out_r_bits_data),
    .io_out_r_bits_last(axi_io_out_r_bits_last),
    .io_icacheio_req(axi_io_icacheio_req),
    .io_icacheio_addr(axi_io_icacheio_addr),
    .io_icacheio_valid(axi_io_icacheio_valid),
    .io_icacheio_data(axi_io_icacheio_data),
    .io_dcacheio_req(axi_io_dcacheio_req),
    .io_dcacheio_raddr(axi_io_dcacheio_raddr),
    .io_dcacheio_rvalid(axi_io_dcacheio_rvalid),
    .io_dcacheio_rdata(axi_io_dcacheio_rdata),
    .io_dcacheio_weq(axi_io_dcacheio_weq),
    .io_dcacheio_waddr(axi_io_dcacheio_waddr),
    .io_dcacheio_wdata(axi_io_dcacheio_wdata),
    .io_dcacheio_wdone(axi_io_dcacheio_wdone)
  );
  Clint clint ( // @[SimTop.scala 20:21]
    .clock(clint_clock),
    .reset(clint_reset),
    .io_dmem_en(clint_io_dmem_en),
    .io_dmem_op(clint_io_dmem_op),
    .io_dmem_addr(clint_io_dmem_addr),
    .io_dmem_wdata(clint_io_dmem_wdata),
    .io_dmem_wmask(clint_io_dmem_wmask),
    .io_dmem_ok(clint_io_dmem_ok),
    .io_dmem_rdata(clint_io_dmem_rdata),
    .io_mem0_en(clint_io_mem0_en),
    .io_mem0_op(clint_io_mem0_op),
    .io_mem0_addr(clint_io_mem0_addr),
    .io_mem0_wdata(clint_io_mem0_wdata),
    .io_mem0_wmask(clint_io_mem0_wmask),
    .io_mem0_ok(clint_io_mem0_ok),
    .io_mem0_rdata(clint_io_mem0_rdata),
    .io_mem1_rdata(clint_io_mem1_rdata),
    .io_mem2_en(clint_io_mem2_en),
    .io_mem2_op(clint_io_mem2_op),
    .io_mem2_wdata(clint_io_mem2_wdata),
    .io_mem2_wmask(clint_io_mem2_wmask),
    .io_mem2_rdata(clint_io_mem2_rdata)
  );
  Mtime mtime ( // @[SimTop.scala 21:21]
    .clock(mtime_clock),
    .reset(mtime_reset),
    .io_mem_rdata(mtime_io_mem_rdata)
  );
  Mtimecmp mtimecmp ( // @[SimTop.scala 22:24]
    .clock(mtimecmp_clock),
    .reset(mtimecmp_reset),
    .io_mem_en(mtimecmp_io_mem_en),
    .io_mem_op(mtimecmp_io_mem_op),
    .io_mem_wdata(mtimecmp_io_mem_wdata),
    .io_mem_wmask(mtimecmp_io_mem_wmask),
    .io_mem_rdata(mtimecmp_io_mem_rdata)
  );
  assign io_uart_out_valid = 1'h0; // @[SimTop.scala 60:21]
  assign io_uart_out_ch = 8'h0; // @[SimTop.scala 61:18]
  assign io_uart_in_valid = 1'h0; // @[SimTop.scala 62:20]
  assign io_memAXI_0_aw_valid = axi_io_out_aw_valid; // @[SimTop.scala 44:17]
  assign io_memAXI_0_aw_bits_len = 8'h7; // @[SimTop.scala 44:17]
  assign io_memAXI_0_aw_bits_size = 3'h3; // @[SimTop.scala 44:17]
  assign io_memAXI_0_aw_bits_burst = 2'h1; // @[SimTop.scala 44:17]
  assign io_memAXI_0_aw_bits_lock = 1'h0; // @[SimTop.scala 44:17]
  assign io_memAXI_0_aw_bits_cache = 4'h2; // @[SimTop.scala 44:17]
  assign io_memAXI_0_aw_bits_qos = 4'h0; // @[SimTop.scala 44:17]
  assign io_memAXI_0_aw_bits_addr = axi_io_out_aw_bits_addr; // @[SimTop.scala 44:17]
  assign io_memAXI_0_aw_bits_prot = 3'h0; // @[SimTop.scala 44:17]
  assign io_memAXI_0_aw_bits_id = 4'h0; // @[SimTop.scala 44:17]
  assign io_memAXI_0_aw_bits_user = 4'h0; // @[SimTop.scala 44:17]
  assign io_memAXI_0_w_valid = axi_io_out_w_valid; // @[SimTop.scala 45:17]
  assign io_memAXI_0_w_bits_data = axi_io_out_w_bits_data; // @[SimTop.scala 45:17]
  assign io_memAXI_0_w_bits_strb = 8'hff; // @[SimTop.scala 45:17]
  assign io_memAXI_0_w_bits_last = axi_io_out_w_bits_last; // @[SimTop.scala 45:17]
  assign io_memAXI_0_b_ready = axi_io_out_b_ready; // @[SimTop.scala 46:17]
  assign io_memAXI_0_ar_valid = axi_io_out_ar_valid; // @[SimTop.scala 42:17]
  assign io_memAXI_0_ar_bits_len = 8'h7; // @[SimTop.scala 42:17]
  assign io_memAXI_0_ar_bits_size = 3'h3; // @[SimTop.scala 42:17]
  assign io_memAXI_0_ar_bits_burst = 2'h1; // @[SimTop.scala 42:17]
  assign io_memAXI_0_ar_bits_lock = 1'h0; // @[SimTop.scala 42:17]
  assign io_memAXI_0_ar_bits_cache = 4'h2; // @[SimTop.scala 42:17]
  assign io_memAXI_0_ar_bits_qos = 4'h0; // @[SimTop.scala 42:17]
  assign io_memAXI_0_ar_bits_addr = axi_io_out_ar_bits_addr; // @[SimTop.scala 42:17]
  assign io_memAXI_0_ar_bits_prot = 3'h0; // @[SimTop.scala 42:17]
  assign io_memAXI_0_ar_bits_id = 4'h0; // @[SimTop.scala 42:17]
  assign io_memAXI_0_ar_bits_user = 4'h0; // @[SimTop.scala 42:17]
  assign io_memAXI_0_r_ready = axi_io_out_r_ready; // @[SimTop.scala 43:17]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_imem_data = icache_io_imem_data; // @[SimTop.scala 26:17]
  assign core_io_imem_data_ok = icache_io_imem_data_ok; // @[SimTop.scala 26:17]
  assign core_io_dmem_ok = clint_io_dmem_ok; // @[SimTop.scala 27:17]
  assign core_io_dmem_rdata = clint_io_dmem_rdata; // @[SimTop.scala 27:17]
  assign icache_clock = clock;
  assign icache_reset = reset;
  assign icache_io_imem_addr = core_io_imem_addr; // @[SimTop.scala 26:17]
  assign icache_io_axi_valid = axi_io_icacheio_valid; // @[SimTop.scala 39:17]
  assign icache_io_axi_data = axi_io_icacheio_data; // @[SimTop.scala 39:17]
  assign dcache_clock = clock;
  assign dcache_reset = reset;
  assign dcache_io_dmem_en = clint_io_mem0_en; // @[SimTop.scala 28:17]
  assign dcache_io_dmem_op = clint_io_mem0_op; // @[SimTop.scala 28:17]
  assign dcache_io_dmem_addr = clint_io_mem0_addr; // @[SimTop.scala 28:17]
  assign dcache_io_dmem_wdata = clint_io_mem0_wdata; // @[SimTop.scala 28:17]
  assign dcache_io_dmem_wmask = clint_io_mem0_wmask; // @[SimTop.scala 28:17]
  assign dcache_io_axi_rvalid = axi_io_dcacheio_rvalid; // @[SimTop.scala 40:17]
  assign dcache_io_axi_rdata = axi_io_dcacheio_rdata; // @[SimTop.scala 40:17]
  assign dcache_io_axi_wdone = axi_io_dcacheio_wdone; // @[SimTop.scala 40:17]
  assign axi_clock = clock;
  assign axi_reset = reset;
  assign axi_io_out_aw_ready = io_memAXI_0_aw_ready; // @[SimTop.scala 44:17]
  assign axi_io_out_w_ready = io_memAXI_0_w_ready; // @[SimTop.scala 45:17]
  assign axi_io_out_b_valid = io_memAXI_0_b_valid; // @[SimTop.scala 46:17]
  assign axi_io_out_ar_ready = io_memAXI_0_ar_ready; // @[SimTop.scala 42:17]
  assign axi_io_out_r_valid = io_memAXI_0_r_valid; // @[SimTop.scala 43:17]
  assign axi_io_out_r_bits_data = io_memAXI_0_r_bits_data; // @[SimTop.scala 43:17]
  assign axi_io_out_r_bits_last = io_memAXI_0_r_bits_last; // @[SimTop.scala 43:17]
  assign axi_io_icacheio_req = icache_io_axi_req; // @[SimTop.scala 39:17]
  assign axi_io_icacheio_addr = icache_io_axi_addr; // @[SimTop.scala 39:17]
  assign axi_io_dcacheio_req = dcache_io_axi_req; // @[SimTop.scala 40:17]
  assign axi_io_dcacheio_raddr = dcache_io_axi_raddr; // @[SimTop.scala 40:17]
  assign axi_io_dcacheio_weq = dcache_io_axi_weq; // @[SimTop.scala 40:17]
  assign axi_io_dcacheio_waddr = dcache_io_axi_waddr; // @[SimTop.scala 40:17]
  assign axi_io_dcacheio_wdata = dcache_io_axi_wdata; // @[SimTop.scala 40:17]
  assign clint_clock = clock;
  assign clint_reset = reset;
  assign clint_io_dmem_en = core_io_dmem_en; // @[SimTop.scala 27:17]
  assign clint_io_dmem_op = core_io_dmem_op; // @[SimTop.scala 27:17]
  assign clint_io_dmem_addr = core_io_dmem_addr; // @[SimTop.scala 27:17]
  assign clint_io_dmem_wdata = core_io_dmem_wdata; // @[SimTop.scala 27:17]
  assign clint_io_dmem_wmask = core_io_dmem_wmask; // @[SimTop.scala 27:17]
  assign clint_io_mem0_ok = dcache_io_dmem_ok; // @[SimTop.scala 28:17]
  assign clint_io_mem0_rdata = dcache_io_dmem_rdata; // @[SimTop.scala 28:17]
  assign clint_io_mem1_rdata = mtime_io_mem_rdata; // @[SimTop.scala 29:17]
  assign clint_io_mem2_rdata = mtimecmp_io_mem_rdata; // @[SimTop.scala 30:17]
  assign mtime_clock = clock;
  assign mtime_reset = reset;
  assign mtimecmp_clock = clock;
  assign mtimecmp_reset = reset;
  assign mtimecmp_io_mem_en = clint_io_mem2_en; // @[SimTop.scala 30:17]
  assign mtimecmp_io_mem_op = clint_io_mem2_op; // @[SimTop.scala 30:17]
  assign mtimecmp_io_mem_wdata = clint_io_mem2_wdata; // @[SimTop.scala 30:17]
  assign mtimecmp_io_mem_wmask = clint_io_mem2_wmask; // @[SimTop.scala 30:17]
endmodule
